// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
neNx+vcxr73XgAY0ToJ43B6ZoS6lf46Lgt8bVZ3IBT63LjI2WNpsr+Co8oACynoGQlsaTswjtKsW
tlVcsM2yAGayMea87+eBsUMO3pYpLFbP90JJk5DFc3OItHz3ttCnb6NSLdah9Xk0rI7w+4RjWaxl
zEHneXmQL+r2ctcsyVuy1eBGzBUWkpD5eIOT/VxfThN7kN+gskpXXmxAvCZW3Lc22bEQqs7HcdFL
ZEe2W5voNJBfluL52A6M32R498y2fkGhYEDhLppL5Z+eIzAgW5ZmoklEodK9KqP1OyWRPh5BHKlI
VsnOsPo3318H7jt/tl/AD2mUwrHoY9Wf5JAl0Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
rU0AVg20scmuYmgT9m+mU2hbdknUqYYkb8itA6rpGOqjoeuYk0fOoNlAovuXEgl6QCWaAfmXo924
aSiDtxPN9blshfe5VQSdFipQV6gO0CZCbLAzCTkuWCrUxHLmRXkImSWLUOdCp/Az+/AltoOTF6m2
xyizuzH4OdfaH5akIEwJZBOoiwnDV1iuWY9Anunrh/1DBEbB4BWShgbeLDNTxJvINTMzs+0tNF0Q
+GRFTuu2/3+Z+Gh+R/ESQYMhihIEJPzALBbGi9VWaGCR68q8/hxyinhDO8b08vmfPVlW7JDLJFQW
EtFQBreZs8ijS+0rjT4bBMFUtT9/Vz0MWpl9+41yFrjSy+PnoJ3LZLwEUuTOQl8An9Cd8scxnAFE
leoDE3HjVzcozUPloYzl6ktOruzVGeOjkoqRscfMJZiaDPXwOfGvrtpL/BJfU01iMLS6EYlV7Soa
ko9l9wJoUeXer3Lrq9PJKNZPDk0d1fAvSLdqBmXQ998cOUp2elH1n2n6fJ/XpoGF/cTqKG0N5u1Q
/HHMLWzfpT3rv/B8hlgai5rNwEOLSrcROpAZt/aHgynssAfn0c9oPT2P4LcsyiVE+wXA1PJxqWqq
FJKb4uYjt66PrzYCw2X8uIW1agLDu8llq6bgrj1ZWbBdws/dDGNvd2VB7GaxM8ip3wwr6eIlVhI8
FBlD6zKjvB6iznSFBKk6hd/E3AOZr5w0wPc0sLgxEC6GgTc9iTwl4+Am7Bfk64J4bzbj2WY0Ntjr
dt40kbAPoXmxq+1c6Y/lK0ks7b1nzWq3gljSK2syfW56ecu6wEbnugM9jkm6WstIfogX1yjAiN78
GSNvYh6zTdwD3Cg1GplfPbz87nySEmwZwvD7fEhIQrGhnfni5w8sCesda985/5qxZnUPgXr+w6hj
XnIk2tPkeBPvqgBgMLlIgpQ2deh2rkGcyF54Uj8hlm11omcnvMhtHVP+J2uN13sJAoLNZy5P3iOD
iERaJEK/WX3vbSXhENSQatj0HZwPN8P46ZwSobSIXbLmwMxfrN17ZqfVVEdkhOVg7mzQ93/O9PCh
1MEVUQCvRrD6Bb1IJptH6+2N9N0FI+zmI9pbV6wzA7u08S3ccYwZL5V/Zix7qxxbZoClOwoZZsDc
dkXOC4lRhsZ8k1VVRM6BfM0uFnygxpd1cMBhA/J/syux7n3nRM+zce3TUqaJcVp00ZkH+ihxV6EE
mMkNK3oCMz7yELpPpgOGMKqRAfkbeeh7sL0HsbiDb79FizBO/ks0S+PEhaupDORXFyfJiNCkvauv
GCo8oME01LWjdnQ1cXGt6jauTxjwzxN/xTiHRLu4BQBfpOS3TgIXjPbRUoNcdOrQjUpTmsKbmnVN
xMTX2SeYsb58bbqwna0YOyr9HiM8Bq9T5MWLYVyXF838SYPo1kvg6jS3LHIqqV1edHskFkJ9e6S1
Fb5eKhbbbsogR0+ygxTVBkPy7yStfIsCUm9sE4n8NM2uuZJTeQ7LkFyPp85BAfh/4RH3Rg6cGovl
ctPKK4TGxwsZHiDGgkRMHRJRZIMsiB8ogqkt2kOiEoh1KQ1ethFXYIIGjshxJW/NCW+DENqVTnYe
Pmww26e50O1tBWh9WhUtFqcQS8gPB4lBHjw+RmxOAOb/xS7sL21q8UttBjfmSiBrTGYTMTvC4puy
5RW+Q3jtis7qoa3gmb+OA7mWWAzXOLsGB5L9Q+d1pnLai2jKhnxqWxl7zg9rG1wECULWSQSm8HVN
1sPB6Tr+z1cstoaSPmSKa8hRwg9BTOtVw+hmwocpPClFDfJhyctS7LzFhsfYlJsppAqMXYzS+SXK
kHJZiO7bBmy54hZakalyaC1vEbb+hMqftlZzQv5XBxefQBOTcnTCwBsjb8csC0sBC2BORj1DSOXI
5TmeqofFxDkLm+fW+clXHBpxzq8dH8U31u2M0RUgqGjBgDr95yIpfhj5oooMMnfIXVNk+I5yLqT9
peZy/eraO4s+JQM1YoSx4L+rNDQN9aPRiPvWkVMCg9XVqlyPIaNPGF4QP1LP3ElhV1niTvkaT8r0
y7Hfwl4jKNkpNpDP9WD8ImJNMLY09Dhv4ZGbTdNU3qeonoNnrEhEElUjkDahzKfpdAYytSFBawtq
QRCylHhT4OohreFJkNGFqwKQDe/e3ICse29SeeD/mp/aEKkww0hW1VJY8dgGupJHKc5TqiBaAtQy
IYk6C+A9jun99g5xwNyywd4AA07CWewUIqHg4d06qWUsVlz7TIpcfzI1bSDUA/wlVYu8BeTbg1mK
QVOzsuHldqeYl3UYD1QBdNb9bIw0AGcZbntgrOynAubRJY5aG0hHtKNwIB1ONu5IstywWVJr9K4D
lWJaauy6AyZWryBUbVdFp0+F3/14LPjE3QlWrxT6Zru1yDb8jqFk49AeAc8sKkgmPIaRNzhUj5QL
lWYP2Wh8FjcpeWAu2kWuL3Is1pTZdUuALLSKhV3dLtciO6M9jhIpgt9r0GbmUvWETndM4D3nGtZJ
uvaakyrXsYoTg1fm0yRqKWzP3KUnv3z2lyGQ9zrcEuwoFJ+NpuXPeqx1sjRpKdjKmVcMyuQ+Uu27
lRrRIItqul4ZmodQ4E32mb0y1mYdWEVFXxVxk4lnF/hWO/gBn1uz9ZftM2Jex+7ii0VY9BYxL1Ni
D8iKjTdReYAZPcn9M4uAln0y321JMk7cKfuwp8byPK4lqODJchEOC0TT0mMh372gb8ulZDC/Y86j
CvbxLzCUv5ah9gDTUwcp9Nd+OYfVv72B9PPIMER8L6SCLbPE68dTHGVVdtzUn/NWH1J5EHmi2aAR
Fc3WI4uYSu9GivhGpbXqlFH8o5WorE/cpWOQ6Yhxu9EXiOoHR7E03TRtUnKU4fOkIzYB0O21ZtEW
6Xf8fZnFDEuTBtzfYbvUmYDZGqTCDUp8W82Yge+5I1xUlhDGtt6c+BgnDqJY7MISBnSx4r6+SWhh
eWvwvjIp6vJTdTlUYu/RePdLHfCODSfp3tdo160XdKgXM5/fjNIQ6saS8lOW+MKqPpyWk6tJbv+C
qb0DUgGGOObI1JkUtYYxWdHfAh3zGULLpxg4OAqIjqhBfaYspTxpwvjEZlQ2LXhLCi5ME+3EgLxT
0/thSepAUjX+ZLg9umlGJbEiB5oYL31A2j+NH0b/HJbY8PTVPmyICzLAvRwRXAhQmdxwu30mYvqZ
rPxlX883S2wU159+u7E5+/u3SoXImKs4yju3jmLEMve4SU3y9c/DfoGCyE5cQNbsMoiFcqIjBWBc
F3QffPNz4emu2xglx9v5X6PDediBHak/0nrOb9d6yS14dgS6avrE+ejpajLukdRjy9KK2g7Qt7KD
59pqG5qlXXxymDycNxP/G4OxGEy6QLT8NmVDcnm9DXjt4diOdHJpxOJUVUO+AYfH4BezDEoeQkjp
wVfw10TQXC35m4U2Gyi/0NAwRMM8VH4AknseGn570mvPm6TDBe4IU8lugj7b9+vvsLktWgUQRISE
wn2cepP7SUrDw5lmlUkWI6FlcweuhEvvyRG5stp99djTlaBEPfJ9BHynRGzLTbsqTCrlcdz8S26f
g+TV5CoVa5p3CoKZMQ8R3hh9OGs+yCPSQvoYTHSPuq9ddO4JxiDHqy4KMeoAhmYa5PeNUOR4mnMa
TWNuJlvBG8SyGNyA1GiLm3awa+DalFun5DqyRb3L//nlnbaOrqb5dCOeO1zC4der9c3ifgAn582T
I8wPNpd5kKXzxRZSG37P9zYJZePV4sHIUaPB8igGxStUxGKCbKBVe6MWLYw1EctzBX94CYmz3EQW
M1kyKNxcDk8wNdvMo+oykVw22wAP2L7tGTYrCUet9Vja5Y/bqp/9/Tc3JgdrR8dEn+6F/KbbmtlN
lnK7EN59sQkN82oKDMK1kCQgVl9rv1DaYwX2NMDjgU8yc8QUI/j8Dph3OknPV/MYX/YpLtLRWKUC
9W4f+lGSusa0KGM7QbvlVZjYDHcM5qtKX2SGzhr5irHs5ZIVLWxEuUy418LVUvbR82rqTfbMXam/
yAAqapsK59GP0tJEInHNAP/KkOBZ2JTRzHFW1dvKVcwBvqf9Lu7pmUnFpTpGlrEllsBKqLoLNWGL
fMfwgIIApP5senoQseZwlQCHCKm7tM7aawFFkgtiJJwT0bcpMaEwd3lYGG9XAPKW/fcLxGZlXtzp
b+SyJRU3th8tVE5D0QnRqtuA1UZIkEpRI/MN2SCfOJBhJkxdd9zOeOahLsm5dCSM53IC/Q+xV3Jz
PHsp729aQOpFu7MuurV4ccthBoHhCVOZYnZRRwhvqKmq3/rcLFM3N/slPkJpja84ZfR6uX9GG0bl
GsBnqJSMHWDUJqlq0/II3hXKqEYsmzNuMwdknbs/1VvLj9gTefH0OirkCTkiET0Gkv3ayozWl+UD
S4u/ocgVDvGePO81slruaszUY2u5HynFfKXQPwOibCpre3wYmzsuKKSBM9NJ/BPsssQfvNMV/AQf
8paHY8NB6k9kIGYjp4WZBRmUvEML+idcPofgnujNtaKhVVq2JTLw7Z770izKdxY/+TR8CtPsSqiT
RT3SYxy/3UOCydWCGX8ER//KJgsOeMyJKlIbgJoOlgCzxJfIuJ9cEqdlWAOqbE9OZzewh/kuv3oN
+kxTvFVhBKtgILzs1JgTDiGKFLGWNs68SEzGyTVfZwSZWF/iIG2v0+LJrdyUoL6+8zH89etYOQ+w
28h/O1nAE1EHuG3QVVaMolTonLxkagIjhP2kR4XTq8BqAf7cC5c2B0V7OUr79Lla+s6DnO8bp8SS
WlFS0Df+7ntxCE9Kn++lmQPyWnP+LrKpizPxT5EcrtPGuMrNc8zsoXq+A2dVkkytNxrcel2JZYqH
VlrUjbxUPuAQDTiqYYYTjH3ZJPdFeTLa2jB53IMVmPUccuwnHhtOVj6Yv6JjNsRgDRZPsAWeLYaW
b4521TvwOtfFpxCQkkBBKavzbzEZ/wWvtkxN1/WML/qZMBtXBhe+cQ+q9DyAEQNTLkxfR1WKXvjc
gspEhCiLZAfZydtjzEPosn79oZh2rgZ9Bocudb8OWHatUsaxmWHFBVn02GyhA7WhJh0JhI4wJzjJ
Rfuw4l9pa/6hxe13RV4aneNMogQXd0ID7p+pUSChdYfBWoNAN2PvQhJmEuhkAG5rGgf5tGye6iNp
ANi/u2GSf49/srqQUprfq7yzTXQm69e95LpBN3Aajs8yOfJR1dj1qNFjsqgNR/bfUO/jNFFyCq9V
kx+00Tb5WNhRoaTckmfr3l5THGstWIKag7yJYb5BDYj/29A2k0umLj/BSwdMR3Bm3pRXYavZw1Nf
zVE756s85ERp8O7dUtDlgryjvYWrYerJ+XkDcfc7IY/qaVRJWZ7pQY3JkYHcmD6YRPcKGu50RCy7
KpkBgi0kmOvKNPatfJVecEiwVr5qfy7MyGf77KnagS7PpV71DkpLDovZebRUMcIxzyWEGeoQpzhK
FUYvvBdhpmcs/9y5x53P0vK0FhL8Lerl0nkhZWRl6u3IjdONy8vAsrNzTg/GsqlDoBIEZBHYf5x8
ZnTQVVVOi2ijJIYBcqRWPtAb3ddBvRtylcKEHNJjfduP2QjY4xLVdEup8YBXwLMp0Xi5B8bHEZRK
XMlAB5+f/wHqLCVOwzeAkoFMkERx3EYyYi6katC1FG1kbOHC/ySd6SwJIF46crNFwbOWrtEdQUYI
LRNSsn4Pmgz60ywnsyz6W4cOjz1qb5WVjv3zFiF0MYwaaOBhtnYcnXn6OhB6F5mov8L2CFvLyUBY
a1rUSEZnUU6n3W3Cs1G09/BVdNYXSdjsH0RgIfIZEujxq9Nv/t/tkKw4VrFcuQHT2pSZxJnY3zP0
betBCsB7gBC/EqCciqkgzJACcBZ+h4ICCZmey/bKYbUb9JEGSEzPyTBhKjILhMAmLVuA3hpRk4Qd
llbFvxamFCJ2IPswga5dP6nO38qvJVKoiJr4/18KCpFFl1iAOC/xRdqrJ2CMWPCbFcn97WNNsO5W
G5YTU0a9fWs1S3SciK1yE2DU+2Ssb9NQqAI01zo7yVWOLfg8oGC54Isvxef4EtEAMDjl2xPP9WdW
kv9rjHrqQi3UZDL7hQlxbfokTC84w/uEuyWFX1gQy9TJJDMEdkZ5Mb1cUVCVPhoOpNViXKFCC6a3
wqrFhoJLXG4Rl0kgzjC9r+u/e+ALfgDIwXkPBI0p/e/t01NuueOseKUl7oUshsR4eS7Ex7QXKd+e
SjUGUPPhRcdq+7dC1dYcmsB2gb0WAXN2MmTH8Nw/nQv2HpgAfxVC32ILNsHoz61iIBxNLvEG4UPj
9IG3HdKN1rsPk5yOtq93jbJNmJByjNVRmXlnoOsoE7gmhqgg+NN5E+UteFtyZXVyiNZI+5MEPcFw
OGbMbsfBQjugy5H/isqSLK9Acw+iQm1+gRR3KnrhGcQdrTt08612RUw8b90EYoR4/Q5SkuEsYzBW
YP/1qlN5fPkDBRC4ToRSuow+nx0KfolX03yJWtlyPz7gKN0uPxUcZLBulrJTQSVJzQh/itWEH+cl
GKDZKPdpOa0k0FBDDQOW8NNN724WhLsJlqE6b4TrKkxsCcL3oq0nt4eH42v+GnE6QzQglU7VThXO
b4uNY5hlyhra2Og82HcYQjV/4L1MJqfQs+3eFSSZZo2Djzk7v7otVd2i6QT7sfXa2pCyRBAx/6ry
0Jpg4U3Loh9dNziJF0o6UXX59gK7LcxRng3PzWU7MlKTs7Vtl7sZsQSLe6wtSavmQxFKll6ewkQi
mdkqYZqxYEnnPt8A3M936AKAgXJ88wjDYTFyVvkSwQ6Jrm3g+40Xz7h3rSSlMcWi9N3M6edANKhI
WK4GmfyKYuaY6/ISwiVxgljKzd7U7fcCfA7sXxzbRioXiA2+9uY905gEU0kGAPBVXYR1/GN+GOZM
MvAA7r3+AUc3pR37GWsvUt8ePY5gnG1AkVrBssKuMlRVH8XaLnxEmSVHg7N5bVzALYhnN6ihETit
grxytINxisrqNFxQCaO1EJQGxVA=
`pragma protect end_protected
