// nios_system.v

// Generated using ACDS version 13.0sp1 232 at 2015.05.23.01:42:12

`timescale 1 ps / 1 ps
module nios_system (
		output wire [6:0]  HEX4_from_the_HEX7_HEX4,                    //       HEX7_HEX4_external_interface.HEX4
		output wire [6:0]  HEX5_from_the_HEX7_HEX4,                    //                                   .HEX5
		output wire [6:0]  HEX6_from_the_HEX7_HEX4,                    //                                   .HEX6
		output wire [6:0]  HEX7_from_the_HEX7_HEX4,                    //                                   .HEX7
		inout  wire [15:0] SRAM_DQ_to_and_from_the_SRAM,               //            SRAM_external_interface.DQ
		output wire [19:0] SRAM_ADDR_from_the_SRAM,                    //                                   .ADDR
		output wire        SRAM_LB_N_from_the_SRAM,                    //                                   .LB_N
		output wire        SRAM_UB_N_from_the_SRAM,                    //                                   .UB_N
		output wire        SRAM_CE_N_from_the_SRAM,                    //                                   .CE_N
		output wire        SRAM_OE_N_from_the_SRAM,                    //                                   .OE_N
		output wire        SRAM_WE_N_from_the_SRAM,                    //                                   .WE_N
		inout  wire [7:0]  LCD_DATA_to_and_from_the_Char_LCD_16x2,     //   Char_LCD_16x2_external_interface.DATA
		output wire        LCD_ON_from_the_Char_LCD_16x2,              //                                   .ON
		output wire        LCD_BLON_from_the_Char_LCD_16x2,            //                                   .BLON
		output wire        LCD_EN_from_the_Char_LCD_16x2,              //                                   .EN
		output wire        LCD_RS_from_the_Char_LCD_16x2,              //                                   .RS
		output wire        LCD_RW_from_the_Char_LCD_16x2,              //                                   .RW
		output wire        sys_clk,                                    //                    sys_clk_out_clk.clk
		input  wire        UART_RXD_to_the_Serial_Port,                //     Serial_Port_external_interface.RXD
		output wire        UART_TXD_from_the_Serial_Port,              //                                   .TXD
		input  wire        AUD_ADCDAT_to_the_Audio,                    //           Audio_external_interface.ADCDAT
		input  wire        AUD_ADCLRCK_to_the_Audio,                   //                                   .ADCLRCK
		input  wire        AUD_BCLK_to_the_Audio,                      //                                   .BCLK
		output wire        AUD_DACDAT_from_the_Audio,                  //                                   .DACDAT
		input  wire        AUD_DACLRCK_to_the_Audio,                   //                                   .DACLRCK
		output wire [17:0] LEDR_from_the_Red_LEDs,                     //        Red_LEDs_external_interface.export
		input  wire        reset_n,                                    //             merged_resets_in_reset.reset_n
		output wire [12:0] zs_addr_from_the_SDRAM,                     //                         SDRAM_wire.addr
		output wire [1:0]  zs_ba_from_the_SDRAM,                       //                                   .ba
		output wire        zs_cas_n_from_the_SDRAM,                    //                                   .cas_n
		output wire        zs_cke_from_the_SDRAM,                      //                                   .cke
		output wire        zs_cs_n_from_the_SDRAM,                     //                                   .cs_n
		inout  wire [31:0] zs_dq_to_and_from_the_SDRAM,                //                                   .dq
		output wire [3:0]  zs_dqm_from_the_SDRAM,                      //                                   .dqm
		output wire        zs_ras_n_from_the_SDRAM,                    //                                   .ras_n
		output wire        zs_we_n_from_the_SDRAM,                     //                                   .we_n
		inout  wire [31:0] GPIO_to_and_from_the_Expansion_JP5,         //   Expansion_JP5_external_interface.export
		output wire [8:0]  LEDG_from_the_Green_LEDs,                   //      Green_LEDs_external_interface.export
		inout  wire        PS2_CLK_to_and_from_the_PS2_Port_Dual,      //   PS2_Port_Dual_external_interface.CLK
		inout  wire        PS2_DAT_to_and_from_the_PS2_Port_Dual,      //                                   .DAT
		input  wire [17:0] Slider_Switches_external_interface_export,  // Slider_Switches_external_interface.export
		inout  wire        I2C_SDAT_to_and_from_the_AV_Config,         //       AV_Config_external_interface.SDAT
		output wire        I2C_SCLK_from_the_AV_Config,                //                                   .SCLK
		inout  wire        PS2_CLK_to_and_from_the_PS2_Port,           //        PS2_Port_external_interface.CLK
		inout  wire        PS2_DAT_to_and_from_the_PS2_Port,           //                                   .DAT
		input  wire [3:0]  KEY_to_the_Pushbuttons,                     //     Pushbuttons_external_interface.export
		input  wire        clk,                                        //                         clk_clk_in.clk
		output wire [6:0]  HEX0_from_the_HEX3_HEX0,                    //       HEX3_HEX0_external_interface.HEX0
		output wire [6:0]  HEX1_from_the_HEX3_HEX0,                    //                                   .HEX1
		output wire [6:0]  HEX2_from_the_HEX3_HEX0,                    //                                   .HEX2
		output wire [6:0]  HEX3_from_the_HEX3_HEX0,                    //                                   .HEX3
		input  wire        clk_27,                                     //                      clk_27_clk_in.clk
		output wire        audio_clk,                                  //                              audio.clk
		output wire        sdram_clk,                                  //                              sdram.clk
		output wire        irda_TXD,                                   //                               irda.TXD
		input  wire        irda_RXD,                                   //                                   .RXD
		inout  wire        sdcard_b_SD_cmd,                            //                             sdcard.b_SD_cmd
		inout  wire        sdcard_b_SD_dat,                            //                                   .b_SD_dat
		inout  wire        sdcard_b_SD_dat3,                           //                                   .b_SD_dat3
		output wire        sdcard_o_SD_clock,                          //                                   .o_SD_clock
		output wire [22:0] flash_ADDR,                                 //                              flash.ADDR
		output wire        flash_CE_N,                                 //                                   .CE_N
		output wire        flash_OE_N,                                 //                                   .OE_N
		output wire        flash_WE_N,                                 //                                   .WE_N
		output wire        flash_RST_N,                                //                                   .RST_N
		inout  wire [7:0]  flash_DQ,                                   //                                   .DQ
		input  wire        video_in_TD_CLK27,                          //                           video_in.TD_CLK27
		input  wire [7:0]  video_in_TD_DATA,                           //                                   .TD_DATA
		input  wire        video_in_TD_HS,                             //                                   .TD_HS
		input  wire        video_in_TD_VS,                             //                                   .TD_VS
		input  wire        video_in_clk27_reset,                       //                                   .clk27_reset
		output wire        video_in_TD_RESET,                          //                                   .TD_RESET
		output wire        video_in_overflow_flag,                     //                                   .overflow_flag
		inout  wire        camera_config_I2C_SDAT,                     //                      camera_config.I2C_SDAT
		output wire        camera_config_I2C_SCLK,                     //                                   .I2C_SCLK
		input  wire [15:0] camera_config_exposure,                     //                                   .exposure
		input  wire        camera_in_PIXEL_CLK,                        //                          camera_in.PIXEL_CLK
		input  wire        camera_in_LINE_VALID,                       //                                   .LINE_VALID
		input  wire        camera_in_FRAME_VALID,                      //                                   .FRAME_VALID
		input  wire        camera_in_pixel_clk_reset,                  //                                   .pixel_clk_reset
		input  wire [11:0] camera_in_PIXEL_DATA,                       //                                   .PIXEL_DATA
		output wire        lcd_controller_external_interface_CLK,      //  lcd_controller_external_interface.CLK
		output wire        lcd_controller_external_interface_HS,       //                                   .HS
		output wire        lcd_controller_external_interface_VS,       //                                   .VS
		output wire        lcd_controller_external_interface_DATA_EN,  //                                   .DATA_EN
		output wire [7:0]  lcd_controller_external_interface_R,        //                                   .R
		output wire [7:0]  lcd_controller_external_interface_G,        //                                   .G
		output wire [7:0]  lcd_controller_external_interface_B,        //                                   .B
		output wire        vga_clk_out_clk_clk,                        //                    vga_clk_out_clk.clk
		inout  wire        accelerometer_I2C_SDAT,                     //                      accelerometer.I2C_SDAT
		output wire        accelerometer_I2C_SCLK,                     //                                   .I2C_SCLK
		output wire        accelerometer_G_SENSOR_CS_N,                //                                   .G_SENSOR_CS_N
		input  wire        accelerometer_G_SENSOR_INT,                 //                                   .G_SENSOR_INT
		input  wire        usb_INT1,                                   //                                usb.INT1
		inout  wire [15:0] usb_DATA,                                   //                                   .DATA
		output wire        usb_RST_N,                                  //                                   .RST_N
		output wire [1:0]  usb_ADDR,                                   //                                   .ADDR
		output wire        usb_CS_N,                                   //                                   .CS_N
		output wire        usb_RD_N,                                   //                                   .RD_N
		output wire        usb_WR_N,                                   //                                   .WR_N
		input  wire        usb_INT0,                                   //                                   .INT0
		output wire        vga_controller_external_interface_CLK,      //  vga_controller_external_interface.CLK
		output wire        vga_controller_external_interface_HS,       //                                   .HS
		output wire        vga_controller_external_interface_VS,       //                                   .VS
		output wire        vga_controller_external_interface_BLANK,    //                                   .BLANK
		output wire        vga_controller_external_interface_SYNC,     //                                   .SYNC
		output wire [7:0]  vga_controller_external_interface_R,        //                                   .R
		output wire [7:0]  vga_controller_external_interface_G,        //                                   .G
		output wire [7:0]  vga_controller_external_interface_B,        //                                   .B
		input  wire        enet_pcs_mac_tx_clk,                        //                    enet_pcs_mac_tx.clk
		input  wire        enet_pcs_mac_rx_clk,                        //                    enet_pcs_mac_rx.clk
		input  wire        enet_mac_status_set_10,                     //                    enet_mac_status.set_10
		input  wire        enet_mac_status_set_1000,                   //                                   .set_1000
		output wire        enet_mac_status_eth_mode,                   //                                   .eth_mode
		output wire        enet_mac_status_ena_10,                     //                                   .ena_10
		input  wire [3:0]  enet_mac_rgmii_rgmii_in,                    //                     enet_mac_rgmii.rgmii_in
		output wire [3:0]  enet_mac_rgmii_rgmii_out,                   //                                   .rgmii_out
		input  wire        enet_mac_rgmii_rx_control,                  //                                   .rx_control
		output wire        enet_mac_rgmii_tx_control,                  //                                   .tx_control
		output wire        enet_mac_mdio_mdc,                          //                      enet_mac_mdio.mdc
		input  wire        enet_mac_mdio_mdio_in,                      //                                   .mdio_in
		output wire        enet_mac_mdio_mdio_out,                     //                                   .mdio_out
		output wire        enet_mac_mdio_mdio_oen,                     //                                   .mdio_oen
		input  wire        enet_mac_misc_xon_gen,                      //                      enet_mac_misc.xon_gen
		input  wire        enet_mac_misc_xoff_gen,                     //                                   .xoff_gen
		output wire        enet_mac_misc_magic_wakeup,                 //                                   .magic_wakeup
		input  wire        enet_mac_misc_magic_sleep_n,                //                                   .magic_sleep_n
		input  wire        enet_mac_misc_ff_tx_crc_fwd,                //                                   .ff_tx_crc_fwd
		output wire        enet_mac_misc_ff_tx_septy,                  //                                   .ff_tx_septy
		output wire        enet_mac_misc_tx_ff_uflow,                  //                                   .tx_ff_uflow
		output wire        enet_mac_misc_ff_tx_a_full,                 //                                   .ff_tx_a_full
		output wire        enet_mac_misc_ff_tx_a_empty,                //                                   .ff_tx_a_empty
		output wire [17:0] enet_mac_misc_rx_err_stat,                  //                                   .rx_err_stat
		output wire [3:0]  enet_mac_misc_rx_frm_type,                  //                                   .rx_frm_type
		output wire        enet_mac_misc_ff_rx_dsav,                   //                                   .ff_rx_dsav
		output wire        enet_mac_misc_ff_rx_a_full,                 //                                   .ff_rx_a_full
		output wire        enet_mac_misc_ff_rx_a_empty,                //                                   .ff_rx_a_empty
		output wire [17:0] videoconferencing_dma_conduit_LEDR_conduit, //      videoconferencing_dma_conduit.LEDR_conduit
		output wire [7:0]  videoconferencing_dma_conduit_LEDG_conduit, //                                   .LEDG_conduit
		output wire [6:0]  videoconferencing_dma_conduit_HEX0_conduit, //                                   .HEX0_conduit
		output wire [6:0]  videoconferencing_dma_conduit_HEX1_conduit, //                                   .HEX1_conduit
		output wire [6:0]  videoconferencing_dma_conduit_HEX2_conduit, //                                   .HEX2_conduit
		output wire [6:0]  videoconferencing_dma_conduit_HEX3_conduit, //                                   .HEX3_conduit
		output wire [6:0]  videoconferencing_dma_conduit_HEX4_conduit, //                                   .HEX4_conduit
		output wire [6:0]  videoconferencing_dma_conduit_HEX5_conduit, //                                   .HEX5_conduit
		output wire [6:0]  videoconferencing_dma_conduit_HEX6_conduit, //                                   .HEX6_conduit
		output wire [6:0]  videoconferencing_dma_conduit_HEX7_conduit, //                                   .HEX7_conduit
		input  wire [17:0] videoconferencing_dma_conduit_SW_conduit    //                                   .SW_conduit
	);

	wire          vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket;                                                                  // VGA_Pixel_RGB_Resampler:stream_out_endofpacket -> VGA_Pixel_Scaler:stream_in_endofpacket
	wire          vga_pixel_rgb_resampler_avalon_rgb_source_valid;                                                                        // VGA_Pixel_RGB_Resampler:stream_out_valid -> VGA_Pixel_Scaler:stream_in_valid
	wire          vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket;                                                                // VGA_Pixel_RGB_Resampler:stream_out_startofpacket -> VGA_Pixel_Scaler:stream_in_startofpacket
	wire   [29:0] vga_pixel_rgb_resampler_avalon_rgb_source_data;                                                                         // VGA_Pixel_RGB_Resampler:stream_out_data -> VGA_Pixel_Scaler:stream_in_data
	wire          vga_pixel_rgb_resampler_avalon_rgb_source_ready;                                                                        // VGA_Pixel_Scaler:stream_in_ready -> VGA_Pixel_RGB_Resampler:stream_out_ready
	wire          vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket;                                                                // VGA_Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	wire          vga_dual_clock_fifo_avalon_dc_buffer_source_valid;                                                                      // VGA_Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	wire          vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket;                                                              // VGA_Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	wire   [29:0] vga_dual_clock_fifo_avalon_dc_buffer_source_data;                                                                       // VGA_Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	wire          vga_dual_clock_fifo_avalon_dc_buffer_source_ready;                                                                      // VGA_Controller:ready -> VGA_Dual_Clock_FIFO:stream_out_ready
	wire          vga_char_buffer_avalon_char_source_endofpacket;                                                                         // VGA_Char_Buffer:stream_endofpacket -> VGA_Alpha_Blender:foreground_endofpacket
	wire          vga_char_buffer_avalon_char_source_valid;                                                                               // VGA_Char_Buffer:stream_valid -> VGA_Alpha_Blender:foreground_valid
	wire          vga_char_buffer_avalon_char_source_startofpacket;                                                                       // VGA_Char_Buffer:stream_startofpacket -> VGA_Alpha_Blender:foreground_startofpacket
	wire   [39:0] vga_char_buffer_avalon_char_source_data;                                                                                // VGA_Char_Buffer:stream_data -> VGA_Alpha_Blender:foreground_data
	wire          vga_char_buffer_avalon_char_source_ready;                                                                               // VGA_Alpha_Blender:foreground_ready -> VGA_Char_Buffer:stream_ready
	wire          vga_pixel_scaler_avalon_scaler_source_endofpacket;                                                                      // VGA_Pixel_Scaler:stream_out_endofpacket -> VGA_Alpha_Blender:background_endofpacket
	wire          vga_pixel_scaler_avalon_scaler_source_valid;                                                                            // VGA_Pixel_Scaler:stream_out_valid -> VGA_Alpha_Blender:background_valid
	wire          vga_pixel_scaler_avalon_scaler_source_startofpacket;                                                                    // VGA_Pixel_Scaler:stream_out_startofpacket -> VGA_Alpha_Blender:background_startofpacket
	wire   [29:0] vga_pixel_scaler_avalon_scaler_source_data;                                                                             // VGA_Pixel_Scaler:stream_out_data -> VGA_Alpha_Blender:background_data
	wire          vga_pixel_scaler_avalon_scaler_source_ready;                                                                            // VGA_Alpha_Blender:background_ready -> VGA_Pixel_Scaler:stream_out_ready
	wire          vga_alpha_blender_avalon_blended_source_endofpacket;                                                                    // VGA_Alpha_Blender:output_endofpacket -> VGA_Dual_Clock_FIFO:stream_in_endofpacket
	wire          vga_alpha_blender_avalon_blended_source_valid;                                                                          // VGA_Alpha_Blender:output_valid -> VGA_Dual_Clock_FIFO:stream_in_valid
	wire          vga_alpha_blender_avalon_blended_source_startofpacket;                                                                  // VGA_Alpha_Blender:output_startofpacket -> VGA_Dual_Clock_FIFO:stream_in_startofpacket
	wire   [29:0] vga_alpha_blender_avalon_blended_source_data;                                                                           // VGA_Alpha_Blender:output_data -> VGA_Dual_Clock_FIFO:stream_in_data
	wire          vga_alpha_blender_avalon_blended_source_ready;                                                                          // VGA_Dual_Clock_FIFO:stream_in_ready -> VGA_Alpha_Blender:output_ready
	wire          video_in_csc_avalon_csc_source_endofpacket;                                                                             // Video_In_CSC:stream_out_endofpacket -> Video_In_RGB_Resampler:stream_in_endofpacket
	wire          video_in_csc_avalon_csc_source_valid;                                                                                   // Video_In_CSC:stream_out_valid -> Video_In_RGB_Resampler:stream_in_valid
	wire          video_in_csc_avalon_csc_source_startofpacket;                                                                           // Video_In_CSC:stream_out_startofpacket -> Video_In_RGB_Resampler:stream_in_startofpacket
	wire   [23:0] video_in_csc_avalon_csc_source_data;                                                                                    // Video_In_CSC:stream_out_data -> Video_In_RGB_Resampler:stream_in_data
	wire          video_in_csc_avalon_csc_source_ready;                                                                                   // Video_In_RGB_Resampler:stream_in_ready -> Video_In_CSC:stream_out_ready
	wire          video_in_rgb_resampler_avalon_rgb_source_endofpacket;                                                                   // Video_In_RGB_Resampler:stream_out_endofpacket -> Video_In_Clipper:stream_in_endofpacket
	wire          video_in_rgb_resampler_avalon_rgb_source_valid;                                                                         // Video_In_RGB_Resampler:stream_out_valid -> Video_In_Clipper:stream_in_valid
	wire          video_in_rgb_resampler_avalon_rgb_source_startofpacket;                                                                 // Video_In_RGB_Resampler:stream_out_startofpacket -> Video_In_Clipper:stream_in_startofpacket
	wire   [15:0] video_in_rgb_resampler_avalon_rgb_source_data;                                                                          // Video_In_RGB_Resampler:stream_out_data -> Video_In_Clipper:stream_in_data
	wire          video_in_rgb_resampler_avalon_rgb_source_ready;                                                                         // Video_In_Clipper:stream_in_ready -> Video_In_RGB_Resampler:stream_out_ready
	wire          video_in_clipper_avalon_clipper_source_endofpacket;                                                                     // Video_In_Clipper:stream_out_endofpacket -> Video_In_Scaler:stream_in_endofpacket
	wire          video_in_clipper_avalon_clipper_source_valid;                                                                           // Video_In_Clipper:stream_out_valid -> Video_In_Scaler:stream_in_valid
	wire          video_in_clipper_avalon_clipper_source_startofpacket;                                                                   // Video_In_Clipper:stream_out_startofpacket -> Video_In_Scaler:stream_in_startofpacket
	wire   [15:0] video_in_clipper_avalon_clipper_source_data;                                                                            // Video_In_Clipper:stream_out_data -> Video_In_Scaler:stream_in_data
	wire          video_in_clipper_avalon_clipper_source_ready;                                                                           // Video_In_Scaler:stream_in_ready -> Video_In_Clipper:stream_out_ready
	wire          video_in_scaler_avalon_scaler_source_endofpacket;                                                                       // Video_In_Scaler:stream_out_endofpacket -> Video_In_DMA_Controller:stream_endofpacket
	wire          video_in_scaler_avalon_scaler_source_valid;                                                                             // Video_In_Scaler:stream_out_valid -> Video_In_DMA_Controller:stream_valid
	wire          video_in_scaler_avalon_scaler_source_startofpacket;                                                                     // Video_In_Scaler:stream_out_startofpacket -> Video_In_DMA_Controller:stream_startofpacket
	wire   [15:0] video_in_scaler_avalon_scaler_source_data;                                                                              // Video_In_Scaler:stream_out_data -> Video_In_DMA_Controller:stream_data
	wire          video_in_scaler_avalon_scaler_source_ready;                                                                             // Video_In_DMA_Controller:stream_ready -> Video_In_Scaler:stream_out_ready
	wire          camera_in_avalon_decoder_source_endofpacket;                                                                            // Camera_In:stream_out_endofpacket -> Camera_Bayer_Resampler:stream_in_endofpacket
	wire          camera_in_avalon_decoder_source_valid;                                                                                  // Camera_In:stream_out_valid -> Camera_Bayer_Resampler:stream_in_valid
	wire          camera_in_avalon_decoder_source_startofpacket;                                                                          // Camera_In:stream_out_startofpacket -> Camera_Bayer_Resampler:stream_in_startofpacket
	wire    [7:0] camera_in_avalon_decoder_source_data;                                                                                   // Camera_In:stream_out_data -> Camera_Bayer_Resampler:stream_in_data
	wire          camera_in_avalon_decoder_source_ready;                                                                                  // Camera_Bayer_Resampler:stream_in_ready -> Camera_In:stream_out_ready
	wire          camera_bayer_resampler_avalon_bayer_source_endofpacket;                                                                 // Camera_Bayer_Resampler:stream_out_endofpacket -> Camera_Scaler:stream_in_endofpacket
	wire          camera_bayer_resampler_avalon_bayer_source_valid;                                                                       // Camera_Bayer_Resampler:stream_out_valid -> Camera_Scaler:stream_in_valid
	wire          camera_bayer_resampler_avalon_bayer_source_startofpacket;                                                               // Camera_Bayer_Resampler:stream_out_startofpacket -> Camera_Scaler:stream_in_startofpacket
	wire   [23:0] camera_bayer_resampler_avalon_bayer_source_data;                                                                        // Camera_Bayer_Resampler:stream_out_data -> Camera_Scaler:stream_in_data
	wire          camera_bayer_resampler_avalon_bayer_source_ready;                                                                       // Camera_Scaler:stream_in_ready -> Camera_Bayer_Resampler:stream_out_ready
	wire          camera_scaler_avalon_scaler_source_endofpacket;                                                                         // Camera_Scaler:stream_out_endofpacket -> Camera_Clipper:stream_in_endofpacket
	wire          camera_scaler_avalon_scaler_source_valid;                                                                               // Camera_Scaler:stream_out_valid -> Camera_Clipper:stream_in_valid
	wire          camera_scaler_avalon_scaler_source_startofpacket;                                                                       // Camera_Scaler:stream_out_startofpacket -> Camera_Clipper:stream_in_startofpacket
	wire   [23:0] camera_scaler_avalon_scaler_source_data;                                                                                // Camera_Scaler:stream_out_data -> Camera_Clipper:stream_in_data
	wire          camera_scaler_avalon_scaler_source_ready;                                                                               // Camera_Clipper:stream_in_ready -> Camera_Scaler:stream_out_ready
	wire          camera_clipper_avalon_clipper_source_endofpacket;                                                                       // Camera_Clipper:stream_out_endofpacket -> Camera_RGB_Resampler:stream_in_endofpacket
	wire          camera_clipper_avalon_clipper_source_valid;                                                                             // Camera_Clipper:stream_out_valid -> Camera_RGB_Resampler:stream_in_valid
	wire          camera_clipper_avalon_clipper_source_startofpacket;                                                                     // Camera_Clipper:stream_out_startofpacket -> Camera_RGB_Resampler:stream_in_startofpacket
	wire   [23:0] camera_clipper_avalon_clipper_source_data;                                                                              // Camera_Clipper:stream_out_data -> Camera_RGB_Resampler:stream_in_data
	wire          camera_clipper_avalon_clipper_source_ready;                                                                             // Camera_RGB_Resampler:stream_in_ready -> Camera_Clipper:stream_out_ready
	wire          camera_rgb_resampler_avalon_rgb_source_endofpacket;                                                                     // Camera_RGB_Resampler:stream_out_endofpacket -> Camera_DMA_Controller:stream_endofpacket
	wire          camera_rgb_resampler_avalon_rgb_source_valid;                                                                           // Camera_RGB_Resampler:stream_out_valid -> Camera_DMA_Controller:stream_valid
	wire          camera_rgb_resampler_avalon_rgb_source_startofpacket;                                                                   // Camera_RGB_Resampler:stream_out_startofpacket -> Camera_DMA_Controller:stream_startofpacket
	wire   [15:0] camera_rgb_resampler_avalon_rgb_source_data;                                                                            // Camera_RGB_Resampler:stream_out_data -> Camera_DMA_Controller:stream_data
	wire          camera_rgb_resampler_avalon_rgb_source_ready;                                                                           // Camera_DMA_Controller:stream_ready -> Camera_RGB_Resampler:stream_out_ready
	wire          external_clocks_vga_clk_33_clk;                                                                                         // External_Clocks:VGA_CLK_33 -> [LCD_Controller:clk, LCD_Dual_Clock_FIFO:clk_stream_out, rst_controller_004:clk]
	wire          lcd_rgb_resampler_avalon_rgb_source_endofpacket;                                                                        // LCD_RGB_Resampler:stream_out_endofpacket -> LCD_Scalar:stream_in_endofpacket
	wire          lcd_rgb_resampler_avalon_rgb_source_valid;                                                                              // LCD_RGB_Resampler:stream_out_valid -> LCD_Scalar:stream_in_valid
	wire          lcd_rgb_resampler_avalon_rgb_source_startofpacket;                                                                      // LCD_RGB_Resampler:stream_out_startofpacket -> LCD_Scalar:stream_in_startofpacket
	wire   [29:0] lcd_rgb_resampler_avalon_rgb_source_data;                                                                               // LCD_RGB_Resampler:stream_out_data -> LCD_Scalar:stream_in_data
	wire          lcd_rgb_resampler_avalon_rgb_source_ready;                                                                              // LCD_Scalar:stream_in_ready -> LCD_RGB_Resampler:stream_out_ready
	wire          lcd_dual_clock_fifo_avalon_dc_buffer_source_endofpacket;                                                                // LCD_Dual_Clock_FIFO:stream_out_endofpacket -> LCD_Controller:endofpacket
	wire          lcd_dual_clock_fifo_avalon_dc_buffer_source_valid;                                                                      // LCD_Dual_Clock_FIFO:stream_out_valid -> LCD_Controller:valid
	wire          lcd_dual_clock_fifo_avalon_dc_buffer_source_startofpacket;                                                              // LCD_Dual_Clock_FIFO:stream_out_startofpacket -> LCD_Controller:startofpacket
	wire   [29:0] lcd_dual_clock_fifo_avalon_dc_buffer_source_data;                                                                       // LCD_Dual_Clock_FIFO:stream_out_data -> LCD_Controller:data
	wire          lcd_dual_clock_fifo_avalon_dc_buffer_source_ready;                                                                      // LCD_Controller:ready -> LCD_Dual_Clock_FIFO:stream_out_ready
	wire          video_in_chroma_resampler_avalon_chroma_source_endofpacket;                                                             // Video_In_Chroma_Resampler:stream_out_endofpacket -> Video_In_CSC:stream_in_endofpacket
	wire          video_in_chroma_resampler_avalon_chroma_source_valid;                                                                   // Video_In_Chroma_Resampler:stream_out_valid -> Video_In_CSC:stream_in_valid
	wire          video_in_chroma_resampler_avalon_chroma_source_startofpacket;                                                           // Video_In_Chroma_Resampler:stream_out_startofpacket -> Video_In_CSC:stream_in_startofpacket
	wire   [23:0] video_in_chroma_resampler_avalon_chroma_source_data;                                                                    // Video_In_Chroma_Resampler:stream_out_data -> Video_In_CSC:stream_in_data
	wire          video_in_chroma_resampler_avalon_chroma_source_ready;                                                                   // Video_In_CSC:stream_in_ready -> Video_In_Chroma_Resampler:stream_out_ready
	wire          video_in_avalon_decoder_source_endofpacket;                                                                             // Video_In:stream_out_endofpacket -> Video_In_Chroma_Resampler:stream_in_endofpacket
	wire          video_in_avalon_decoder_source_valid;                                                                                   // Video_In:stream_out_valid -> Video_In_Chroma_Resampler:stream_in_valid
	wire          video_in_avalon_decoder_source_startofpacket;                                                                           // Video_In:stream_out_startofpacket -> Video_In_Chroma_Resampler:stream_in_startofpacket
	wire   [15:0] video_in_avalon_decoder_source_data;                                                                                    // Video_In:stream_out_data -> Video_In_Chroma_Resampler:stream_in_data
	wire          video_in_avalon_decoder_source_ready;                                                                                   // Video_In_Chroma_Resampler:stream_in_ready -> Video_In:stream_out_ready
	wire          lcd_alpha_blender_avalon_blended_source_endofpacket;                                                                    // LCD_Alpha_Blender:output_endofpacket -> LCD_Dual_Clock_FIFO:stream_in_endofpacket
	wire          lcd_alpha_blender_avalon_blended_source_valid;                                                                          // LCD_Alpha_Blender:output_valid -> LCD_Dual_Clock_FIFO:stream_in_valid
	wire          lcd_alpha_blender_avalon_blended_source_startofpacket;                                                                  // LCD_Alpha_Blender:output_startofpacket -> LCD_Dual_Clock_FIFO:stream_in_startofpacket
	wire   [29:0] lcd_alpha_blender_avalon_blended_source_data;                                                                           // LCD_Alpha_Blender:output_data -> LCD_Dual_Clock_FIFO:stream_in_data
	wire          lcd_alpha_blender_avalon_blended_source_ready;                                                                          // LCD_Dual_Clock_FIFO:stream_in_ready -> LCD_Alpha_Blender:output_ready
	wire          lcd_scalar_avalon_scaler_source_endofpacket;                                                                            // LCD_Scalar:stream_out_endofpacket -> LCD_Alpha_Blender:background_endofpacket
	wire          lcd_scalar_avalon_scaler_source_valid;                                                                                  // LCD_Scalar:stream_out_valid -> LCD_Alpha_Blender:background_valid
	wire          lcd_scalar_avalon_scaler_source_startofpacket;                                                                          // LCD_Scalar:stream_out_startofpacket -> LCD_Alpha_Blender:background_startofpacket
	wire   [29:0] lcd_scalar_avalon_scaler_source_data;                                                                                   // LCD_Scalar:stream_out_data -> LCD_Alpha_Blender:background_data
	wire          lcd_scalar_avalon_scaler_source_ready;                                                                                  // LCD_Alpha_Blender:background_ready -> LCD_Scalar:stream_out_ready
	wire          lcd_char_buffer_avalon_char_source_endofpacket;                                                                         // LCD_Char_Buffer:stream_endofpacket -> LCD_Alpha_Blender:foreground_endofpacket
	wire          lcd_char_buffer_avalon_char_source_valid;                                                                               // LCD_Char_Buffer:stream_valid -> LCD_Alpha_Blender:foreground_valid
	wire          lcd_char_buffer_avalon_char_source_startofpacket;                                                                       // LCD_Char_Buffer:stream_startofpacket -> LCD_Alpha_Blender:foreground_startofpacket
	wire   [39:0] lcd_char_buffer_avalon_char_source_data;                                                                                // LCD_Char_Buffer:stream_data -> LCD_Alpha_Blender:foreground_data
	wire          lcd_char_buffer_avalon_char_source_ready;                                                                               // LCD_Alpha_Blender:foreground_ready -> LCD_Char_Buffer:stream_ready
	wire          cpu_jtag_debug_module_reset_reset;                                                                                      // CPU:jtag_debug_module_resetrequest -> [LCD_DMA_Controller:reset, LCD_DMA_Controller_avalon_dma_control_slave_translator:reset, LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:reset, LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LCD_DMA_Controller_avalon_dma_master_translator:reset, LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:reset, VGA_DMA_Controller:reset, VGA_DMA_Controller_avalon_dma_control_slave_translator:reset, VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:reset, VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_DMA_Controller_avalon_dma_master_translator:reset, VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:reset, addr_router_004:reset, addr_router_005:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, id_router_035:reset, id_router_036:reset, rsp_xbar_demux_035:reset, rsp_xbar_demux_036:reset, rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in3, rst_controller_003:reset_in1, rst_controller_004:reset_in1, rst_controller_005:reset_in1]
	wire          lcd_dma_controller_avalon_pixel_source_endofpacket;                                                                     // LCD_DMA_Controller:stream_endofpacket -> LCD_RGB_Resampler:stream_in_endofpacket
	wire          lcd_dma_controller_avalon_pixel_source_valid;                                                                           // LCD_DMA_Controller:stream_valid -> LCD_RGB_Resampler:stream_in_valid
	wire          lcd_dma_controller_avalon_pixel_source_startofpacket;                                                                   // LCD_DMA_Controller:stream_startofpacket -> LCD_RGB_Resampler:stream_in_startofpacket
	wire   [15:0] lcd_dma_controller_avalon_pixel_source_data;                                                                            // LCD_DMA_Controller:stream_data -> LCD_RGB_Resampler:stream_in_data
	wire          lcd_dma_controller_avalon_pixel_source_ready;                                                                           // LCD_RGB_Resampler:stream_in_ready -> LCD_DMA_Controller:stream_ready
	wire          vga_dma_controller_avalon_pixel_source_endofpacket;                                                                     // VGA_DMA_Controller:stream_endofpacket -> VGA_Pixel_RGB_Resampler:stream_in_endofpacket
	wire          vga_dma_controller_avalon_pixel_source_valid;                                                                           // VGA_DMA_Controller:stream_valid -> VGA_Pixel_RGB_Resampler:stream_in_valid
	wire          vga_dma_controller_avalon_pixel_source_startofpacket;                                                                   // VGA_DMA_Controller:stream_startofpacket -> VGA_Pixel_RGB_Resampler:stream_in_startofpacket
	wire   [15:0] vga_dma_controller_avalon_pixel_source_data;                                                                            // VGA_DMA_Controller:stream_data -> VGA_Pixel_RGB_Resampler:stream_in_data
	wire          vga_dma_controller_avalon_pixel_source_ready;                                                                           // VGA_Pixel_RGB_Resampler:stream_in_ready -> VGA_DMA_Controller:stream_ready
	wire          cpu_custom_instruction_master_multi_readra;                                                                             // CPU:A_ci_multi_readra -> CPU_custom_instruction_master_translator:ci_slave_multi_readra
	wire    [7:0] cpu_custom_instruction_master_multi_n;                                                                                  // CPU:A_ci_multi_n -> CPU_custom_instruction_master_translator:ci_slave_multi_n
	wire          cpu_custom_instruction_master_multi_readrb;                                                                             // CPU:A_ci_multi_readrb -> CPU_custom_instruction_master_translator:ci_slave_multi_readrb
	wire          cpu_custom_instruction_master_done;                                                                                     // CPU_custom_instruction_master_translator:ci_slave_multi_done -> CPU:A_ci_multi_done
	wire          cpu_custom_instruction_master_clk_en;                                                                                   // CPU:A_ci_multi_clk_en -> CPU_custom_instruction_master_translator:ci_slave_multi_clken
	wire          cpu_custom_instruction_master_multi_writerc;                                                                            // CPU:A_ci_multi_writerc -> CPU_custom_instruction_master_translator:ci_slave_multi_writerc
	wire   [31:0] cpu_custom_instruction_master_multi_result;                                                                             // CPU_custom_instruction_master_translator:ci_slave_multi_result -> CPU:A_ci_multi_result
	wire          cpu_custom_instruction_master_clk;                                                                                      // CPU:A_ci_multi_clock -> CPU_custom_instruction_master_translator:ci_slave_multi_clk
	wire    [4:0] cpu_custom_instruction_master_multi_c;                                                                                  // CPU:A_ci_multi_c -> CPU_custom_instruction_master_translator:ci_slave_multi_c
	wire    [4:0] cpu_custom_instruction_master_multi_b;                                                                                  // CPU:A_ci_multi_b -> CPU_custom_instruction_master_translator:ci_slave_multi_b
	wire    [4:0] cpu_custom_instruction_master_multi_a;                                                                                  // CPU:A_ci_multi_a -> CPU_custom_instruction_master_translator:ci_slave_multi_a
	wire   [31:0] cpu_custom_instruction_master_multi_dataa;                                                                              // CPU:A_ci_multi_dataa -> CPU_custom_instruction_master_translator:ci_slave_multi_dataa
	wire          cpu_custom_instruction_master_start;                                                                                    // CPU:A_ci_multi_start -> CPU_custom_instruction_master_translator:ci_slave_multi_start
	wire   [31:0] cpu_custom_instruction_master_multi_datab;                                                                              // CPU:A_ci_multi_datab -> CPU_custom_instruction_master_translator:ci_slave_multi_datab
	wire          cpu_custom_instruction_master_reset;                                                                                    // CPU:A_ci_multi_reset -> CPU_custom_instruction_master_translator:ci_slave_multi_reset
	wire   [31:0] cpu_custom_instruction_master_translator_multi_ci_master_result;                                                        // CPU_custom_instruction_master_multi_xconnect:ci_slave_result -> CPU_custom_instruction_master_translator:multi_ci_master_result
	wire    [4:0] cpu_custom_instruction_master_translator_multi_ci_master_b;                                                             // CPU_custom_instruction_master_translator:multi_ci_master_b -> CPU_custom_instruction_master_multi_xconnect:ci_slave_b
	wire    [4:0] cpu_custom_instruction_master_translator_multi_ci_master_c;                                                             // CPU_custom_instruction_master_translator:multi_ci_master_c -> CPU_custom_instruction_master_multi_xconnect:ci_slave_c
	wire          cpu_custom_instruction_master_translator_multi_ci_master_clk_en;                                                        // CPU_custom_instruction_master_translator:multi_ci_master_clken -> CPU_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire          cpu_custom_instruction_master_translator_multi_ci_master_done;                                                          // CPU_custom_instruction_master_multi_xconnect:ci_slave_done -> CPU_custom_instruction_master_translator:multi_ci_master_done
	wire    [4:0] cpu_custom_instruction_master_translator_multi_ci_master_a;                                                             // CPU_custom_instruction_master_translator:multi_ci_master_a -> CPU_custom_instruction_master_multi_xconnect:ci_slave_a
	wire    [7:0] cpu_custom_instruction_master_translator_multi_ci_master_n;                                                             // CPU_custom_instruction_master_translator:multi_ci_master_n -> CPU_custom_instruction_master_multi_xconnect:ci_slave_n
	wire          cpu_custom_instruction_master_translator_multi_ci_master_writerc;                                                       // CPU_custom_instruction_master_translator:multi_ci_master_writerc -> CPU_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire          cpu_custom_instruction_master_translator_multi_ci_master_clk;                                                           // CPU_custom_instruction_master_translator:multi_ci_master_clk -> CPU_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire          cpu_custom_instruction_master_translator_multi_ci_master_start;                                                         // CPU_custom_instruction_master_translator:multi_ci_master_start -> CPU_custom_instruction_master_multi_xconnect:ci_slave_start
	wire   [31:0] cpu_custom_instruction_master_translator_multi_ci_master_dataa;                                                         // CPU_custom_instruction_master_translator:multi_ci_master_dataa -> CPU_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire          cpu_custom_instruction_master_translator_multi_ci_master_readra;                                                        // CPU_custom_instruction_master_translator:multi_ci_master_readra -> CPU_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire          cpu_custom_instruction_master_translator_multi_ci_master_reset;                                                         // CPU_custom_instruction_master_translator:multi_ci_master_reset -> CPU_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire   [31:0] cpu_custom_instruction_master_translator_multi_ci_master_datab;                                                         // CPU_custom_instruction_master_translator:multi_ci_master_datab -> CPU_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire          cpu_custom_instruction_master_translator_multi_ci_master_readrb;                                                        // CPU_custom_instruction_master_translator:multi_ci_master_readrb -> CPU_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_result;                                                         // CPU_custom_instruction_master_multi_slave_translator0:ci_slave_result -> CPU_custom_instruction_master_multi_xconnect:ci_master0_result
	wire    [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_b;                                                              // CPU_custom_instruction_master_multi_xconnect:ci_master0_b -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire    [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_c;                                                              // CPU_custom_instruction_master_multi_xconnect:ci_master0_c -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire          cpu_custom_instruction_master_multi_xconnect_ci_master0_done;                                                           // CPU_custom_instruction_master_multi_slave_translator0:ci_slave_done -> CPU_custom_instruction_master_multi_xconnect:ci_master0_done
	wire          cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en;                                                         // CPU_custom_instruction_master_multi_xconnect:ci_master0_clken -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire    [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_a;                                                              // CPU_custom_instruction_master_multi_xconnect:ci_master0_a -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire    [7:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_n;                                                              // CPU_custom_instruction_master_multi_xconnect:ci_master0_n -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire          cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc;                                                        // CPU_custom_instruction_master_multi_xconnect:ci_master0_writerc -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire   [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending;                                                       // CPU_custom_instruction_master_multi_xconnect:ci_master0_ipending -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire          cpu_custom_instruction_master_multi_xconnect_ci_master0_clk;                                                            // CPU_custom_instruction_master_multi_xconnect:ci_master0_clk -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire          cpu_custom_instruction_master_multi_xconnect_ci_master0_start;                                                          // CPU_custom_instruction_master_multi_xconnect:ci_master0_start -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire   [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa;                                                          // CPU_custom_instruction_master_multi_xconnect:ci_master0_dataa -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire          cpu_custom_instruction_master_multi_xconnect_ci_master0_readra;                                                         // CPU_custom_instruction_master_multi_xconnect:ci_master0_readra -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire          cpu_custom_instruction_master_multi_xconnect_ci_master0_reset;                                                          // CPU_custom_instruction_master_multi_xconnect:ci_master0_reset -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire   [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_datab;                                                          // CPU_custom_instruction_master_multi_xconnect:ci_master0_datab -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire          cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb;                                                         // CPU_custom_instruction_master_multi_xconnect:ci_master0_readrb -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire          cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus;                                                        // CPU_custom_instruction_master_multi_xconnect:ci_master0_estatus -> CPU_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire   [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_result;                                                 // CPU_fpoint:result -> CPU_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire          cpu_custom_instruction_master_multi_slave_translator0_ci_master_start;                                                  // CPU_custom_instruction_master_multi_slave_translator0:ci_master_start -> CPU_fpoint:start
	wire   [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa;                                                  // CPU_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> CPU_fpoint:dataa
	wire          cpu_custom_instruction_master_multi_slave_translator0_ci_master_done;                                                   // CPU_fpoint:done -> CPU_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire          cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;                                                 // CPU_custom_instruction_master_multi_slave_translator0:ci_master_clken -> CPU_fpoint:clk_en
	wire    [1:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_n;                                                      // CPU_custom_instruction_master_multi_slave_translator0:ci_master_n -> CPU_fpoint:n
	wire          cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset;                                                  // CPU_custom_instruction_master_multi_slave_translator0:ci_master_reset -> CPU_fpoint:reset
	wire   [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab;                                                  // CPU_custom_instruction_master_multi_slave_translator0:ci_master_datab -> CPU_fpoint:datab
	wire          cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk;                                                    // CPU_custom_instruction_master_multi_slave_translator0:ci_master_clk -> CPU_fpoint:clk
	wire          cpu_instruction_master_waitrequest;                                                                                     // CPU_instruction_master_translator:av_waitrequest -> CPU:i_waitrequest
	wire   [27:0] cpu_instruction_master_address;                                                                                         // CPU:i_address -> CPU_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                                            // CPU:i_read -> CPU_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                                        // CPU_instruction_master_translator:av_readdata -> CPU:i_readdata
	wire          cpu_instruction_master_readdatavalid;                                                                                   // CPU_instruction_master_translator:av_readdatavalid -> CPU:i_readdatavalid
	wire          cpu_data_master_waitrequest;                                                                                            // CPU_data_master_translator:av_waitrequest -> CPU:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                                              // CPU:d_writedata -> CPU_data_master_translator:av_writedata
	wire   [28:0] cpu_data_master_address;                                                                                                // CPU:d_address -> CPU_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                                                  // CPU:d_write -> CPU_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                                                   // CPU:d_read -> CPU_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                                               // CPU_data_master_translator:av_readdata -> CPU:d_readdata
	wire          cpu_data_master_debugaccess;                                                                                            // CPU:jtag_debug_module_debugaccess_to_roms -> CPU_data_master_translator:av_debugaccess
	wire    [3:0] cpu_data_master_byteenable;                                                                                             // CPU:d_byteenable -> CPU_data_master_translator:av_byteenable
	wire          video_in_dma_controller_avalon_dma_master_waitrequest;                                                                  // Video_In_DMA_Controller_avalon_dma_master_translator:av_waitrequest -> Video_In_DMA_Controller:master_waitrequest
	wire   [15:0] video_in_dma_controller_avalon_dma_master_writedata;                                                                    // Video_In_DMA_Controller:master_writedata -> Video_In_DMA_Controller_avalon_dma_master_translator:av_writedata
	wire   [31:0] video_in_dma_controller_avalon_dma_master_address;                                                                      // Video_In_DMA_Controller:master_address -> Video_In_DMA_Controller_avalon_dma_master_translator:av_address
	wire          video_in_dma_controller_avalon_dma_master_write;                                                                        // Video_In_DMA_Controller:master_write -> Video_In_DMA_Controller_avalon_dma_master_translator:av_write
	wire          camera_dma_controller_avalon_dma_master_waitrequest;                                                                    // Camera_DMA_Controller_avalon_dma_master_translator:av_waitrequest -> Camera_DMA_Controller:master_waitrequest
	wire   [15:0] camera_dma_controller_avalon_dma_master_writedata;                                                                      // Camera_DMA_Controller:master_writedata -> Camera_DMA_Controller_avalon_dma_master_translator:av_writedata
	wire   [31:0] camera_dma_controller_avalon_dma_master_address;                                                                        // Camera_DMA_Controller:master_address -> Camera_DMA_Controller_avalon_dma_master_translator:av_address
	wire          camera_dma_controller_avalon_dma_master_write;                                                                          // Camera_DMA_Controller:master_write -> Camera_DMA_Controller_avalon_dma_master_translator:av_write
	wire          lcd_dma_controller_avalon_dma_master_waitrequest;                                                                       // LCD_DMA_Controller_avalon_dma_master_translator:av_waitrequest -> LCD_DMA_Controller:master_waitrequest
	wire   [31:0] lcd_dma_controller_avalon_dma_master_address;                                                                           // LCD_DMA_Controller:master_address -> LCD_DMA_Controller_avalon_dma_master_translator:av_address
	wire          lcd_dma_controller_avalon_dma_master_lock;                                                                              // LCD_DMA_Controller:master_arbiterlock -> LCD_DMA_Controller_avalon_dma_master_translator:av_lock
	wire          lcd_dma_controller_avalon_dma_master_read;                                                                              // LCD_DMA_Controller:master_read -> LCD_DMA_Controller_avalon_dma_master_translator:av_read
	wire   [15:0] lcd_dma_controller_avalon_dma_master_readdata;                                                                          // LCD_DMA_Controller_avalon_dma_master_translator:av_readdata -> LCD_DMA_Controller:master_readdata
	wire          lcd_dma_controller_avalon_dma_master_readdatavalid;                                                                     // LCD_DMA_Controller_avalon_dma_master_translator:av_readdatavalid -> LCD_DMA_Controller:master_readdatavalid
	wire          vga_dma_controller_avalon_dma_master_waitrequest;                                                                       // VGA_DMA_Controller_avalon_dma_master_translator:av_waitrequest -> VGA_DMA_Controller:master_waitrequest
	wire   [31:0] vga_dma_controller_avalon_dma_master_address;                                                                           // VGA_DMA_Controller:master_address -> VGA_DMA_Controller_avalon_dma_master_translator:av_address
	wire          vga_dma_controller_avalon_dma_master_lock;                                                                              // VGA_DMA_Controller:master_arbiterlock -> VGA_DMA_Controller_avalon_dma_master_translator:av_lock
	wire          vga_dma_controller_avalon_dma_master_read;                                                                              // VGA_DMA_Controller:master_read -> VGA_DMA_Controller_avalon_dma_master_translator:av_read
	wire   [15:0] vga_dma_controller_avalon_dma_master_readdata;                                                                          // VGA_DMA_Controller_avalon_dma_master_translator:av_readdata -> VGA_DMA_Controller:master_readdata
	wire          vga_dma_controller_avalon_dma_master_readdatavalid;                                                                     // VGA_DMA_Controller_avalon_dma_master_translator:av_readdatavalid -> VGA_DMA_Controller:master_readdatavalid
	wire          videoconferencing_dma_0_avalon_master_waitrequest;                                                                      // VideoConferencing_DMA_0_avalon_master_translator:av_waitrequest -> VideoConferencing_DMA_0:master_waitrequest
	wire   [15:0] videoconferencing_dma_0_avalon_master_writedata;                                                                        // VideoConferencing_DMA_0:master_writedata -> VideoConferencing_DMA_0_avalon_master_translator:av_writedata
	wire   [31:0] videoconferencing_dma_0_avalon_master_address;                                                                          // VideoConferencing_DMA_0:master_address -> VideoConferencing_DMA_0_avalon_master_translator:av_address
	wire          videoconferencing_dma_0_avalon_master_write;                                                                            // VideoConferencing_DMA_0:master_write -> VideoConferencing_DMA_0_avalon_master_translator:av_write
	wire    [1:0] videoconferencing_dma_0_avalon_master_byteenable;                                                                       // VideoConferencing_DMA_0:master_byteenable -> VideoConferencing_DMA_0_avalon_master_translator:av_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                                       // CPU:jtag_debug_module_waitrequest -> CPU_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                                         // CPU_jtag_debug_module_translator:av_writedata -> CPU:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                                           // CPU_jtag_debug_module_translator:av_address -> CPU:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                             // CPU_jtag_debug_module_translator:av_write -> CPU:jtag_debug_module_write
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_read;                                                              // CPU_jtag_debug_module_translator:av_read -> CPU:jtag_debug_module_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                                          // CPU:jtag_debug_module_readdata -> CPU_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                                       // CPU_jtag_debug_module_translator:av_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                                        // CPU_jtag_debug_module_translator:av_byteenable -> CPU:jtag_debug_module_byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                                    // SDRAM:za_waitrequest -> SDRAM_s1_translator:av_waitrequest
	wire   [31:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                                      // SDRAM_s1_translator:av_writedata -> SDRAM:az_data
	wire   [24:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                                        // SDRAM_s1_translator:av_address -> SDRAM:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                                     // SDRAM_s1_translator:av_chipselect -> SDRAM:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                                          // SDRAM_s1_translator:av_write -> SDRAM:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                                           // SDRAM_s1_translator:av_read -> SDRAM:az_rd_n
	wire   [31:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                                       // SDRAM:za_data -> SDRAM_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                                  // SDRAM:za_valid -> SDRAM_s1_translator:av_readdatavalid
	wire    [3:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                                     // SDRAM_s1_translator:av_byteenable -> SDRAM:az_be_n
	wire          flash_flash_data_translator_avalon_anti_slave_0_waitrequest;                                                            // Flash:o_avalon_waitrequest -> Flash_flash_data_translator:av_waitrequest
	wire   [31:0] flash_flash_data_translator_avalon_anti_slave_0_writedata;                                                              // Flash_flash_data_translator:av_writedata -> Flash:i_avalon_writedata
	wire   [20:0] flash_flash_data_translator_avalon_anti_slave_0_address;                                                                // Flash_flash_data_translator:av_address -> Flash:i_avalon_address
	wire          flash_flash_data_translator_avalon_anti_slave_0_chipselect;                                                             // Flash_flash_data_translator:av_chipselect -> Flash:i_avalon_chip_select
	wire          flash_flash_data_translator_avalon_anti_slave_0_write;                                                                  // Flash_flash_data_translator:av_write -> Flash:i_avalon_write
	wire          flash_flash_data_translator_avalon_anti_slave_0_read;                                                                   // Flash_flash_data_translator:av_read -> Flash:i_avalon_read
	wire   [31:0] flash_flash_data_translator_avalon_anti_slave_0_readdata;                                                               // Flash:o_avalon_readdata -> Flash_flash_data_translator:av_readdata
	wire    [3:0] flash_flash_data_translator_avalon_anti_slave_0_byteenable;                                                             // Flash_flash_data_translator:av_byteenable -> Flash:i_avalon_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                                 // JTAG_UART:av_waitrequest -> JTAG_UART_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                                   // JTAG_UART_avalon_jtag_slave_translator:av_writedata -> JTAG_UART:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                                     // JTAG_UART_avalon_jtag_slave_translator:av_address -> JTAG_UART:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                                  // JTAG_UART_avalon_jtag_slave_translator:av_chipselect -> JTAG_UART:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                                       // JTAG_UART_avalon_jtag_slave_translator:av_write -> JTAG_UART:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                                        // JTAG_UART_avalon_jtag_slave_translator:av_read -> JTAG_UART:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                                    // JTAG_UART:av_readdata -> JTAG_UART_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] interval_timer_s1_translator_avalon_anti_slave_0_writedata;                                                             // Interval_Timer_s1_translator:av_writedata -> Interval_Timer:writedata
	wire    [2:0] interval_timer_s1_translator_avalon_anti_slave_0_address;                                                               // Interval_Timer_s1_translator:av_address -> Interval_Timer:address
	wire          interval_timer_s1_translator_avalon_anti_slave_0_chipselect;                                                            // Interval_Timer_s1_translator:av_chipselect -> Interval_Timer:chipselect
	wire          interval_timer_s1_translator_avalon_anti_slave_0_write;                                                                 // Interval_Timer_s1_translator:av_write -> Interval_Timer:write_n
	wire   [15:0] interval_timer_s1_translator_avalon_anti_slave_0_readdata;                                                              // Interval_Timer:readdata -> Interval_Timer_s1_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                                             // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                                            // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [31:0] red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                           // Red_LEDs_avalon_parallel_port_slave_translator:av_writedata -> Red_LEDs:writedata
	wire    [1:0] red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                             // Red_LEDs_avalon_parallel_port_slave_translator:av_address -> Red_LEDs:address
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                          // Red_LEDs_avalon_parallel_port_slave_translator:av_chipselect -> Red_LEDs:chipselect
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                               // Red_LEDs_avalon_parallel_port_slave_translator:av_write -> Red_LEDs:write
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                                // Red_LEDs_avalon_parallel_port_slave_translator:av_read -> Red_LEDs:read
	wire   [31:0] red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                            // Red_LEDs:readdata -> Red_LEDs_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                          // Red_LEDs_avalon_parallel_port_slave_translator:av_byteenable -> Red_LEDs:byteenable
	wire   [31:0] green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                         // Green_LEDs_avalon_parallel_port_slave_translator:av_writedata -> Green_LEDs:writedata
	wire    [1:0] green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                           // Green_LEDs_avalon_parallel_port_slave_translator:av_address -> Green_LEDs:address
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                        // Green_LEDs_avalon_parallel_port_slave_translator:av_chipselect -> Green_LEDs:chipselect
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                             // Green_LEDs_avalon_parallel_port_slave_translator:av_write -> Green_LEDs:write
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                              // Green_LEDs_avalon_parallel_port_slave_translator:av_read -> Green_LEDs:read
	wire   [31:0] green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                          // Green_LEDs:readdata -> Green_LEDs_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                        // Green_LEDs_avalon_parallel_port_slave_translator:av_byteenable -> Green_LEDs:byteenable
	wire   [31:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                          // HEX3_HEX0_avalon_parallel_port_slave_translator:av_writedata -> HEX3_HEX0:writedata
	wire    [1:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                            // HEX3_HEX0_avalon_parallel_port_slave_translator:av_address -> HEX3_HEX0:address
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                         // HEX3_HEX0_avalon_parallel_port_slave_translator:av_chipselect -> HEX3_HEX0:chipselect
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                              // HEX3_HEX0_avalon_parallel_port_slave_translator:av_write -> HEX3_HEX0:write
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                               // HEX3_HEX0_avalon_parallel_port_slave_translator:av_read -> HEX3_HEX0:read
	wire   [31:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                           // HEX3_HEX0:readdata -> HEX3_HEX0_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                         // HEX3_HEX0_avalon_parallel_port_slave_translator:av_byteenable -> HEX3_HEX0:byteenable
	wire   [31:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                          // HEX7_HEX4_avalon_parallel_port_slave_translator:av_writedata -> HEX7_HEX4:writedata
	wire    [1:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                            // HEX7_HEX4_avalon_parallel_port_slave_translator:av_address -> HEX7_HEX4:address
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                         // HEX7_HEX4_avalon_parallel_port_slave_translator:av_chipselect -> HEX7_HEX4:chipselect
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                              // HEX7_HEX4_avalon_parallel_port_slave_translator:av_write -> HEX7_HEX4:write
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                               // HEX7_HEX4_avalon_parallel_port_slave_translator:av_read -> HEX7_HEX4:read
	wire   [31:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                           // HEX7_HEX4:readdata -> HEX7_HEX4_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                         // HEX7_HEX4_avalon_parallel_port_slave_translator:av_byteenable -> HEX7_HEX4:byteenable
	wire   [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                    // Slider_Switches_avalon_parallel_port_slave_translator:av_writedata -> Slider_Switches:writedata
	wire    [1:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                      // Slider_Switches_avalon_parallel_port_slave_translator:av_address -> Slider_Switches:address
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                   // Slider_Switches_avalon_parallel_port_slave_translator:av_chipselect -> Slider_Switches:chipselect
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                        // Slider_Switches_avalon_parallel_port_slave_translator:av_write -> Slider_Switches:write
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                         // Slider_Switches_avalon_parallel_port_slave_translator:av_read -> Slider_Switches:read
	wire   [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                     // Slider_Switches:readdata -> Slider_Switches_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                   // Slider_Switches_avalon_parallel_port_slave_translator:av_byteenable -> Slider_Switches:byteenable
	wire   [31:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                        // Pushbuttons_avalon_parallel_port_slave_translator:av_writedata -> Pushbuttons:writedata
	wire    [1:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                          // Pushbuttons_avalon_parallel_port_slave_translator:av_address -> Pushbuttons:address
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                       // Pushbuttons_avalon_parallel_port_slave_translator:av_chipselect -> Pushbuttons:chipselect
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                            // Pushbuttons_avalon_parallel_port_slave_translator:av_write -> Pushbuttons:write
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                             // Pushbuttons_avalon_parallel_port_slave_translator:av_read -> Pushbuttons:read
	wire   [31:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                         // Pushbuttons:readdata -> Pushbuttons_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                       // Pushbuttons_avalon_parallel_port_slave_translator:av_byteenable -> Pushbuttons:byteenable
	wire   [31:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata;                                      // Expansion_JP5_avalon_parallel_port_slave_translator:av_writedata -> Expansion_JP5:writedata
	wire    [1:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address;                                        // Expansion_JP5_avalon_parallel_port_slave_translator:av_address -> Expansion_JP5:address
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect;                                     // Expansion_JP5_avalon_parallel_port_slave_translator:av_chipselect -> Expansion_JP5:chipselect
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write;                                          // Expansion_JP5_avalon_parallel_port_slave_translator:av_write -> Expansion_JP5:write
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read;                                           // Expansion_JP5_avalon_parallel_port_slave_translator:av_read -> Expansion_JP5:read
	wire   [31:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata;                                       // Expansion_JP5:readdata -> Expansion_JP5_avalon_parallel_port_slave_translator:av_readdata
	wire    [3:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable;                                     // Expansion_JP5_avalon_parallel_port_slave_translator:av_byteenable -> Expansion_JP5:byteenable
	wire   [31:0] serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata;                                                // Serial_Port_avalon_rs232_slave_translator:av_writedata -> Serial_Port:writedata
	wire    [0:0] serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_address;                                                  // Serial_Port_avalon_rs232_slave_translator:av_address -> Serial_Port:address
	wire          serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect;                                               // Serial_Port_avalon_rs232_slave_translator:av_chipselect -> Serial_Port:chipselect
	wire          serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_write;                                                    // Serial_Port_avalon_rs232_slave_translator:av_write -> Serial_Port:write
	wire          serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_read;                                                     // Serial_Port_avalon_rs232_slave_translator:av_read -> Serial_Port:read
	wire   [31:0] serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata;                                                 // Serial_Port:readdata -> Serial_Port_avalon_rs232_slave_translator:av_readdata
	wire    [3:0] serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable;                                               // Serial_Port_avalon_rs232_slave_translator:av_byteenable -> Serial_Port:byteenable
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest;                                              // Char_LCD_16x2:waitrequest -> Char_LCD_16x2_avalon_lcd_slave_translator:av_waitrequest
	wire    [7:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata;                                                // Char_LCD_16x2_avalon_lcd_slave_translator:av_writedata -> Char_LCD_16x2:writedata
	wire    [0:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_address;                                                  // Char_LCD_16x2_avalon_lcd_slave_translator:av_address -> Char_LCD_16x2:address
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect;                                               // Char_LCD_16x2_avalon_lcd_slave_translator:av_chipselect -> Char_LCD_16x2:chipselect
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_write;                                                    // Char_LCD_16x2_avalon_lcd_slave_translator:av_write -> Char_LCD_16x2:write
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_read;                                                     // Char_LCD_16x2_avalon_lcd_slave_translator:av_read -> Char_LCD_16x2:read
	wire    [7:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata;                                                 // Char_LCD_16x2:readdata -> Char_LCD_16x2_avalon_lcd_slave_translator:av_readdata
	wire          ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest;                                                   // PS2_Port:waitrequest -> PS2_Port_avalon_ps2_slave_translator:av_waitrequest
	wire   [31:0] ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata;                                                     // PS2_Port_avalon_ps2_slave_translator:av_writedata -> PS2_Port:writedata
	wire    [0:0] ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_address;                                                       // PS2_Port_avalon_ps2_slave_translator:av_address -> PS2_Port:address
	wire          ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect;                                                    // PS2_Port_avalon_ps2_slave_translator:av_chipselect -> PS2_Port:chipselect
	wire          ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_write;                                                         // PS2_Port_avalon_ps2_slave_translator:av_write -> PS2_Port:write
	wire          ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_read;                                                          // PS2_Port_avalon_ps2_slave_translator:av_read -> PS2_Port:read
	wire   [31:0] ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata;                                                      // PS2_Port:readdata -> PS2_Port_avalon_ps2_slave_translator:av_readdata
	wire    [3:0] ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable;                                                    // PS2_Port_avalon_ps2_slave_translator:av_byteenable -> PS2_Port:byteenable
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                                        // SRAM_avalon_sram_slave_translator:av_writedata -> SRAM:writedata
	wire   [19:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                                          // SRAM_avalon_sram_slave_translator:av_address -> SRAM:address
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                                            // SRAM_avalon_sram_slave_translator:av_write -> SRAM:write
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                                             // SRAM_avalon_sram_slave_translator:av_read -> SRAM:read
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                                         // SRAM:readdata -> SRAM_avalon_sram_slave_translator:av_readdata
	wire          sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                                    // SRAM:readdatavalid -> SRAM_avalon_sram_slave_translator:av_readdatavalid
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                                       // SRAM_avalon_sram_slave_translator:av_byteenable -> SRAM:byteenable
	wire   [31:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata;                                     // VGA_Char_Buffer_avalon_char_control_slave_translator:av_writedata -> VGA_Char_Buffer:ctrl_writedata
	wire    [0:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address;                                       // VGA_Char_Buffer_avalon_char_control_slave_translator:av_address -> VGA_Char_Buffer:ctrl_address
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect;                                    // VGA_Char_Buffer_avalon_char_control_slave_translator:av_chipselect -> VGA_Char_Buffer:ctrl_chipselect
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write;                                         // VGA_Char_Buffer_avalon_char_control_slave_translator:av_write -> VGA_Char_Buffer:ctrl_write
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read;                                          // VGA_Char_Buffer_avalon_char_control_slave_translator:av_read -> VGA_Char_Buffer:ctrl_read
	wire   [31:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata;                                      // VGA_Char_Buffer:ctrl_readdata -> VGA_Char_Buffer_avalon_char_control_slave_translator:av_readdata
	wire    [3:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable;                                    // VGA_Char_Buffer_avalon_char_control_slave_translator:av_byteenable -> VGA_Char_Buffer:ctrl_byteenable
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest;                                    // VGA_Char_Buffer:buf_waitrequest -> VGA_Char_Buffer_avalon_char_buffer_slave_translator:av_waitrequest
	wire    [7:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata;                                      // VGA_Char_Buffer_avalon_char_buffer_slave_translator:av_writedata -> VGA_Char_Buffer:buf_writedata
	wire   [12:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address;                                        // VGA_Char_Buffer_avalon_char_buffer_slave_translator:av_address -> VGA_Char_Buffer:buf_address
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect;                                     // VGA_Char_Buffer_avalon_char_buffer_slave_translator:av_chipselect -> VGA_Char_Buffer:buf_chipselect
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write;                                          // VGA_Char_Buffer_avalon_char_buffer_slave_translator:av_write -> VGA_Char_Buffer:buf_write
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read;                                           // VGA_Char_Buffer_avalon_char_buffer_slave_translator:av_read -> VGA_Char_Buffer:buf_read
	wire    [7:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata;                                       // VGA_Char_Buffer:buf_readdata -> VGA_Char_Buffer_avalon_char_buffer_slave_translator:av_readdata
	wire    [0:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable;                                     // VGA_Char_Buffer_avalon_char_buffer_slave_translator:av_byteenable -> VGA_Char_Buffer:buf_byteenable
	wire          onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest;                                           // OnBoard_AV:waitrequest -> OnBoard_AV_avalon_av_config_slave_translator:av_waitrequest
	wire   [31:0] onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata;                                             // OnBoard_AV_avalon_av_config_slave_translator:av_writedata -> OnBoard_AV:writedata
	wire    [1:0] onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_address;                                               // OnBoard_AV_avalon_av_config_slave_translator:av_address -> OnBoard_AV:address
	wire          onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_write;                                                 // OnBoard_AV_avalon_av_config_slave_translator:av_write -> OnBoard_AV:write
	wire          onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_read;                                                  // OnBoard_AV_avalon_av_config_slave_translator:av_read -> OnBoard_AV:read
	wire   [31:0] onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata;                                              // OnBoard_AV:readdata -> OnBoard_AV_avalon_av_config_slave_translator:av_readdata
	wire    [3:0] onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable;                                            // OnBoard_AV_avalon_av_config_slave_translator:av_byteenable -> OnBoard_AV:byteenable
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest;                                              // PS2_Port_Dual:waitrequest -> PS2_Port_Dual_avalon_ps2_slave_translator:av_waitrequest
	wire   [31:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata;                                                // PS2_Port_Dual_avalon_ps2_slave_translator:av_writedata -> PS2_Port_Dual:writedata
	wire    [0:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_address;                                                  // PS2_Port_Dual_avalon_ps2_slave_translator:av_address -> PS2_Port_Dual:address
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect;                                               // PS2_Port_Dual_avalon_ps2_slave_translator:av_chipselect -> PS2_Port_Dual:chipselect
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_write;                                                    // PS2_Port_Dual_avalon_ps2_slave_translator:av_write -> PS2_Port_Dual:write
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_read;                                                     // PS2_Port_Dual_avalon_ps2_slave_translator:av_read -> PS2_Port_Dual:read
	wire   [31:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata;                                                 // PS2_Port_Dual:readdata -> PS2_Port_Dual_avalon_ps2_slave_translator:av_readdata
	wire    [3:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable;                                               // PS2_Port_Dual_avalon_ps2_slave_translator:av_byteenable -> PS2_Port_Dual:byteenable
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_anti_slave_0_writedata;                                                      // Audio_avalon_audio_slave_translator:av_writedata -> Audio:writedata
	wire    [1:0] audio_avalon_audio_slave_translator_avalon_anti_slave_0_address;                                                        // Audio_avalon_audio_slave_translator:av_address -> Audio:address
	wire          audio_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect;                                                     // Audio_avalon_audio_slave_translator:av_chipselect -> Audio:chipselect
	wire          audio_avalon_audio_slave_translator_avalon_anti_slave_0_write;                                                          // Audio_avalon_audio_slave_translator:av_write -> Audio:write
	wire          audio_avalon_audio_slave_translator_avalon_anti_slave_0_read;                                                           // Audio_avalon_audio_slave_translator:av_read -> Audio:read
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_anti_slave_0_readdata;                                                       // Audio:readdata -> Audio_avalon_audio_slave_translator:av_readdata
	wire          flash_flash_erase_control_translator_avalon_anti_slave_0_waitrequest;                                                   // Flash:o_avalon_erase_waitrequest -> Flash_flash_erase_control_translator:av_waitrequest
	wire   [31:0] flash_flash_erase_control_translator_avalon_anti_slave_0_writedata;                                                     // Flash_flash_erase_control_translator:av_writedata -> Flash:i_avalon_erase_writedata
	wire          flash_flash_erase_control_translator_avalon_anti_slave_0_chipselect;                                                    // Flash_flash_erase_control_translator:av_chipselect -> Flash:i_avalon_erase_chip_select
	wire          flash_flash_erase_control_translator_avalon_anti_slave_0_write;                                                         // Flash_flash_erase_control_translator:av_write -> Flash:i_avalon_erase_write
	wire          flash_flash_erase_control_translator_avalon_anti_slave_0_read;                                                          // Flash_flash_erase_control_translator:av_read -> Flash:i_avalon_erase_read
	wire   [31:0] flash_flash_erase_control_translator_avalon_anti_slave_0_readdata;                                                      // Flash:o_avalon_erase_readdata -> Flash_flash_erase_control_translator:av_readdata
	wire    [3:0] flash_flash_erase_control_translator_avalon_anti_slave_0_byteenable;                                                    // Flash_flash_erase_control_translator:av_byteenable -> Flash:i_avalon_erase_byteenable
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest;                                                 // SD_Card:o_avalon_waitrequest -> SD_Card_avalon_sdcard_slave_translator:av_waitrequest
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata;                                                   // SD_Card_avalon_sdcard_slave_translator:av_writedata -> SD_Card:i_avalon_writedata
	wire    [7:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address;                                                     // SD_Card_avalon_sdcard_slave_translator:av_address -> SD_Card:i_avalon_address
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect;                                                  // SD_Card_avalon_sdcard_slave_translator:av_chipselect -> SD_Card:i_avalon_chip_select
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write;                                                       // SD_Card_avalon_sdcard_slave_translator:av_write -> SD_Card:i_avalon_write
	wire          sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read;                                                        // SD_Card_avalon_sdcard_slave_translator:av_read -> SD_Card:i_avalon_read
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata;                                                    // SD_Card:o_avalon_readdata -> SD_Card_avalon_sdcard_slave_translator:av_readdata
	wire    [3:0] sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable;                                                  // SD_Card_avalon_sdcard_slave_translator:av_byteenable -> SD_Card:i_avalon_byteenable
	wire   [31:0] irda_avalon_irda_slave_translator_avalon_anti_slave_0_writedata;                                                        // IrDA_avalon_irda_slave_translator:av_writedata -> IrDA:writedata
	wire    [0:0] irda_avalon_irda_slave_translator_avalon_anti_slave_0_address;                                                          // IrDA_avalon_irda_slave_translator:av_address -> IrDA:address
	wire          irda_avalon_irda_slave_translator_avalon_anti_slave_0_chipselect;                                                       // IrDA_avalon_irda_slave_translator:av_chipselect -> IrDA:chipselect
	wire          irda_avalon_irda_slave_translator_avalon_anti_slave_0_write;                                                            // IrDA_avalon_irda_slave_translator:av_write -> IrDA:write
	wire          irda_avalon_irda_slave_translator_avalon_anti_slave_0_read;                                                             // IrDA_avalon_irda_slave_translator:av_read -> IrDA:read
	wire   [31:0] irda_avalon_irda_slave_translator_avalon_anti_slave_0_readdata;                                                         // IrDA:readdata -> IrDA_avalon_irda_slave_translator:av_readdata
	wire    [3:0] irda_avalon_irda_slave_translator_avalon_anti_slave_0_byteenable;                                                       // IrDA_avalon_irda_slave_translator:av_byteenable -> IrDA:byteenable
	wire   [31:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata;                              // Video_In_DMA_Controller_avalon_dma_control_slave_translator:av_writedata -> Video_In_DMA_Controller:slave_writedata
	wire    [1:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address;                                // Video_In_DMA_Controller_avalon_dma_control_slave_translator:av_address -> Video_In_DMA_Controller:slave_address
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write;                                  // Video_In_DMA_Controller_avalon_dma_control_slave_translator:av_write -> Video_In_DMA_Controller:slave_write
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read;                                   // Video_In_DMA_Controller_avalon_dma_control_slave_translator:av_read -> Video_In_DMA_Controller:slave_read
	wire   [31:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata;                               // Video_In_DMA_Controller:slave_readdata -> Video_In_DMA_Controller_avalon_dma_control_slave_translator:av_readdata
	wire    [3:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable;                             // Video_In_DMA_Controller_avalon_dma_control_slave_translator:av_byteenable -> Video_In_DMA_Controller:slave_byteenable
	wire   [31:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata;                                // Camera_DMA_Controller_avalon_dma_control_slave_translator:av_writedata -> Camera_DMA_Controller:slave_writedata
	wire    [1:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address;                                  // Camera_DMA_Controller_avalon_dma_control_slave_translator:av_address -> Camera_DMA_Controller:slave_address
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write;                                    // Camera_DMA_Controller_avalon_dma_control_slave_translator:av_write -> Camera_DMA_Controller:slave_write
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read;                                     // Camera_DMA_Controller_avalon_dma_control_slave_translator:av_read -> Camera_DMA_Controller:slave_read
	wire   [31:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata;                                 // Camera_DMA_Controller:slave_readdata -> Camera_DMA_Controller_avalon_dma_control_slave_translator:av_readdata
	wire    [3:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable;                               // Camera_DMA_Controller_avalon_dma_control_slave_translator:av_byteenable -> Camera_DMA_Controller:slave_byteenable
	wire          camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest;                                        // Camera_Config:waitrequest -> Camera_Config_avalon_av_config_slave_translator:av_waitrequest
	wire   [31:0] camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata;                                          // Camera_Config_avalon_av_config_slave_translator:av_writedata -> Camera_Config:writedata
	wire    [1:0] camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address;                                            // Camera_Config_avalon_av_config_slave_translator:av_address -> Camera_Config:address
	wire          camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write;                                              // Camera_Config_avalon_av_config_slave_translator:av_write -> Camera_Config:write
	wire          camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read;                                               // Camera_Config_avalon_av_config_slave_translator:av_read -> Camera_Config:read
	wire   [31:0] camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata;                                           // Camera_Config:readdata -> Camera_Config_avalon_av_config_slave_translator:av_readdata
	wire    [3:0] camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable;                                         // Camera_Config_avalon_av_config_slave_translator:av_byteenable -> Camera_Config:byteenable
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_waitrequest;                           // Accelerometer:waitrequest -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator:av_waitrequest
	wire    [7:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_writedata;                             // Accelerometer_avalon_accelerometer_spi_mode_slave_translator:av_writedata -> Accelerometer:writedata
	wire    [0:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_address;                               // Accelerometer_avalon_accelerometer_spi_mode_slave_translator:av_address -> Accelerometer:address
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_write;                                 // Accelerometer_avalon_accelerometer_spi_mode_slave_translator:av_write -> Accelerometer:write
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_read;                                  // Accelerometer_avalon_accelerometer_spi_mode_slave_translator:av_read -> Accelerometer:read
	wire    [7:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_readdata;                              // Accelerometer:readdata -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator:av_readdata
	wire    [0:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_byteenable;                            // Accelerometer_avalon_accelerometer_spi_mode_slave_translator:av_byteenable -> Accelerometer:byteenable
	wire   [15:0] usb_avalon_usb_slave_translator_avalon_anti_slave_0_writedata;                                                          // USB_avalon_usb_slave_translator:av_writedata -> USB:writedata
	wire    [1:0] usb_avalon_usb_slave_translator_avalon_anti_slave_0_address;                                                            // USB_avalon_usb_slave_translator:av_address -> USB:address
	wire          usb_avalon_usb_slave_translator_avalon_anti_slave_0_chipselect;                                                         // USB_avalon_usb_slave_translator:av_chipselect -> USB:chipselect
	wire          usb_avalon_usb_slave_translator_avalon_anti_slave_0_write;                                                              // USB_avalon_usb_slave_translator:av_write -> USB:write
	wire          usb_avalon_usb_slave_translator_avalon_anti_slave_0_read;                                                               // USB_avalon_usb_slave_translator:av_read -> USB:read
	wire   [15:0] usb_avalon_usb_slave_translator_avalon_anti_slave_0_readdata;                                                           // USB:readdata -> USB_avalon_usb_slave_translator:av_readdata
	wire   [31:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata;                                     // LCD_Char_Buffer_avalon_char_control_slave_translator:av_writedata -> LCD_Char_Buffer:ctrl_writedata
	wire    [0:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address;                                       // LCD_Char_Buffer_avalon_char_control_slave_translator:av_address -> LCD_Char_Buffer:ctrl_address
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect;                                    // LCD_Char_Buffer_avalon_char_control_slave_translator:av_chipselect -> LCD_Char_Buffer:ctrl_chipselect
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write;                                         // LCD_Char_Buffer_avalon_char_control_slave_translator:av_write -> LCD_Char_Buffer:ctrl_write
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read;                                          // LCD_Char_Buffer_avalon_char_control_slave_translator:av_read -> LCD_Char_Buffer:ctrl_read
	wire   [31:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata;                                      // LCD_Char_Buffer:ctrl_readdata -> LCD_Char_Buffer_avalon_char_control_slave_translator:av_readdata
	wire    [3:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable;                                    // LCD_Char_Buffer_avalon_char_control_slave_translator:av_byteenable -> LCD_Char_Buffer:ctrl_byteenable
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest;                                    // LCD_Char_Buffer:buf_waitrequest -> LCD_Char_Buffer_avalon_char_buffer_slave_translator:av_waitrequest
	wire    [7:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata;                                      // LCD_Char_Buffer_avalon_char_buffer_slave_translator:av_writedata -> LCD_Char_Buffer:buf_writedata
	wire   [10:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address;                                        // LCD_Char_Buffer_avalon_char_buffer_slave_translator:av_address -> LCD_Char_Buffer:buf_address
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect;                                     // LCD_Char_Buffer_avalon_char_buffer_slave_translator:av_chipselect -> LCD_Char_Buffer:buf_chipselect
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write;                                          // LCD_Char_Buffer_avalon_char_buffer_slave_translator:av_write -> LCD_Char_Buffer:buf_write
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read;                                           // LCD_Char_Buffer_avalon_char_buffer_slave_translator:av_read -> LCD_Char_Buffer:buf_read
	wire    [7:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata;                                       // LCD_Char_Buffer:buf_readdata -> LCD_Char_Buffer_avalon_char_buffer_slave_translator:av_readdata
	wire    [0:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable;                                     // LCD_Char_Buffer_avalon_char_buffer_slave_translator:av_byteenable -> LCD_Char_Buffer:buf_byteenable
	wire          enet_control_port_translator_avalon_anti_slave_0_waitrequest;                                                           // enet:waitrequest -> enet_control_port_translator:av_waitrequest
	wire   [31:0] enet_control_port_translator_avalon_anti_slave_0_writedata;                                                             // enet_control_port_translator:av_writedata -> enet:writedata
	wire    [7:0] enet_control_port_translator_avalon_anti_slave_0_address;                                                               // enet_control_port_translator:av_address -> enet:address
	wire          enet_control_port_translator_avalon_anti_slave_0_write;                                                                 // enet_control_port_translator:av_write -> enet:write
	wire          enet_control_port_translator_avalon_anti_slave_0_read;                                                                  // enet_control_port_translator:av_read -> enet:read
	wire   [31:0] enet_control_port_translator_avalon_anti_slave_0_readdata;                                                              // enet:readdata -> enet_control_port_translator:av_readdata
	wire   [31:0] packet_memory_s1_translator_avalon_anti_slave_0_writedata;                                                              // packet_memory_s1_translator:av_writedata -> packet_memory:writedata
	wire    [9:0] packet_memory_s1_translator_avalon_anti_slave_0_address;                                                                // packet_memory_s1_translator:av_address -> packet_memory:address
	wire          packet_memory_s1_translator_avalon_anti_slave_0_chipselect;                                                             // packet_memory_s1_translator:av_chipselect -> packet_memory:chipselect
	wire          packet_memory_s1_translator_avalon_anti_slave_0_clken;                                                                  // packet_memory_s1_translator:av_clken -> packet_memory:clken
	wire          packet_memory_s1_translator_avalon_anti_slave_0_write;                                                                  // packet_memory_s1_translator:av_write -> packet_memory:write
	wire   [31:0] packet_memory_s1_translator_avalon_anti_slave_0_readdata;                                                               // packet_memory:readdata -> packet_memory_s1_translator:av_readdata
	wire    [3:0] packet_memory_s1_translator_avalon_anti_slave_0_byteenable;                                                             // packet_memory_s1_translator:av_byteenable -> packet_memory:byteenable
	wire   [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_writedata;                                                          // descriptor_memory_s1_translator:av_writedata -> descriptor_memory:writedata
	wire    [9:0] descriptor_memory_s1_translator_avalon_anti_slave_0_address;                                                            // descriptor_memory_s1_translator:av_address -> descriptor_memory:address
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect;                                                         // descriptor_memory_s1_translator:av_chipselect -> descriptor_memory:chipselect
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_clken;                                                              // descriptor_memory_s1_translator:av_clken -> descriptor_memory:clken
	wire          descriptor_memory_s1_translator_avalon_anti_slave_0_write;                                                              // descriptor_memory_s1_translator:av_write -> descriptor_memory:write
	wire   [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_readdata;                                                           // descriptor_memory:readdata -> descriptor_memory_s1_translator:av_readdata
	wire    [3:0] descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable;                                                         // descriptor_memory_s1_translator:av_byteenable -> descriptor_memory:byteenable
	wire   [31:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata;                                   // LCD_DMA_Controller_avalon_dma_control_slave_translator:av_writedata -> LCD_DMA_Controller:slave_writedata
	wire    [1:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address;                                     // LCD_DMA_Controller_avalon_dma_control_slave_translator:av_address -> LCD_DMA_Controller:slave_address
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write;                                       // LCD_DMA_Controller_avalon_dma_control_slave_translator:av_write -> LCD_DMA_Controller:slave_write
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read;                                        // LCD_DMA_Controller_avalon_dma_control_slave_translator:av_read -> LCD_DMA_Controller:slave_read
	wire   [31:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata;                                    // LCD_DMA_Controller:slave_readdata -> LCD_DMA_Controller_avalon_dma_control_slave_translator:av_readdata
	wire    [3:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable;                                  // LCD_DMA_Controller_avalon_dma_control_slave_translator:av_byteenable -> LCD_DMA_Controller:slave_byteenable
	wire   [31:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata;                                   // VGA_DMA_Controller_avalon_dma_control_slave_translator:av_writedata -> VGA_DMA_Controller:slave_writedata
	wire    [1:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address;                                     // VGA_DMA_Controller_avalon_dma_control_slave_translator:av_address -> VGA_DMA_Controller:slave_address
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write;                                       // VGA_DMA_Controller_avalon_dma_control_slave_translator:av_write -> VGA_DMA_Controller:slave_write
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read;                                        // VGA_DMA_Controller_avalon_dma_control_slave_translator:av_read -> VGA_DMA_Controller:slave_read
	wire   [31:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata;                                    // VGA_DMA_Controller:slave_readdata -> VGA_DMA_Controller_avalon_dma_control_slave_translator:av_readdata
	wire    [3:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable;                                  // VGA_DMA_Controller_avalon_dma_control_slave_translator:av_byteenable -> VGA_DMA_Controller:slave_byteenable
	wire   [31:0] videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_writedata;                                          // VideoConferencing_DMA_0_avalon_slave_translator:av_writedata -> VideoConferencing_DMA_0:slave_writedata
	wire    [7:0] videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_address;                                            // VideoConferencing_DMA_0_avalon_slave_translator:av_address -> VideoConferencing_DMA_0:slave_address
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_chipselect;                                         // VideoConferencing_DMA_0_avalon_slave_translator:av_chipselect -> VideoConferencing_DMA_0:slave_chipselect
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_write;                                              // VideoConferencing_DMA_0_avalon_slave_translator:av_write -> VideoConferencing_DMA_0:slave_write
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_read;                                               // VideoConferencing_DMA_0_avalon_slave_translator:av_read -> VideoConferencing_DMA_0:slave_read
	wire   [31:0] videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_readdata;                                           // VideoConferencing_DMA_0:slave_readdata -> VideoConferencing_DMA_0_avalon_slave_translator:av_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                                                // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                                                 // CPU_instruction_master_translator:uav_burstcount -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                                                  // CPU_instruction_master_translator:uav_writedata -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                                    // CPU_instruction_master_translator:uav_address -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                                       // CPU_instruction_master_translator:uav_lock -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                                      // CPU_instruction_master_translator:uav_write -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                                       // CPU_instruction_master_translator:uav_read -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                                                   // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                                                // CPU_instruction_master_translator:uav_debugaccess -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                                                 // CPU_instruction_master_translator:uav_byteenable -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                              // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_instruction_master_translator:uav_readdatavalid
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                                       // CPU_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                                        // CPU_data_master_translator:uav_burstcount -> CPU_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                                         // CPU_data_master_translator:uav_writedata -> CPU_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_address;                                                           // CPU_data_master_translator:uav_address -> CPU_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                                              // CPU_data_master_translator:uav_lock -> CPU_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                                             // CPU_data_master_translator:uav_write -> CPU_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                                              // CPU_data_master_translator:uav_read -> CPU_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                                          // CPU_data_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                                       // CPU_data_master_translator:uav_debugaccess -> CPU_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                                        // CPU_data_master_translator:uav_byteenable -> CPU_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                                     // CPU_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_data_master_translator:uav_readdatavalid
	wire          video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest;                             // Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> Video_In_DMA_Controller_avalon_dma_master_translator:uav_waitrequest
	wire    [1:0] video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount;                              // Video_In_DMA_Controller_avalon_dma_master_translator:uav_burstcount -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata;                               // Video_In_DMA_Controller_avalon_dma_master_translator:uav_writedata -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address;                                 // Video_In_DMA_Controller_avalon_dma_master_translator:uav_address -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock;                                    // Video_In_DMA_Controller_avalon_dma_master_translator:uav_lock -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write;                                   // Video_In_DMA_Controller_avalon_dma_master_translator:uav_write -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read;                                    // Video_In_DMA_Controller_avalon_dma_master_translator:uav_read -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata;                                // Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> Video_In_DMA_Controller_avalon_dma_master_translator:uav_readdata
	wire          video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess;                             // Video_In_DMA_Controller_avalon_dma_master_translator:uav_debugaccess -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable;                              // Video_In_DMA_Controller_avalon_dma_master_translator:uav_byteenable -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid;                           // Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> Video_In_DMA_Controller_avalon_dma_master_translator:uav_readdatavalid
	wire          camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest;                               // Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> Camera_DMA_Controller_avalon_dma_master_translator:uav_waitrequest
	wire    [1:0] camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount;                                // Camera_DMA_Controller_avalon_dma_master_translator:uav_burstcount -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata;                                 // Camera_DMA_Controller_avalon_dma_master_translator:uav_writedata -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address;                                   // Camera_DMA_Controller_avalon_dma_master_translator:uav_address -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock;                                      // Camera_DMA_Controller_avalon_dma_master_translator:uav_lock -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write;                                     // Camera_DMA_Controller_avalon_dma_master_translator:uav_write -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read;                                      // Camera_DMA_Controller_avalon_dma_master_translator:uav_read -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata;                                  // Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> Camera_DMA_Controller_avalon_dma_master_translator:uav_readdata
	wire          camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess;                               // Camera_DMA_Controller_avalon_dma_master_translator:uav_debugaccess -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable;                                // Camera_DMA_Controller_avalon_dma_master_translator:uav_byteenable -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid;                             // Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> Camera_DMA_Controller_avalon_dma_master_translator:uav_readdatavalid
	wire          lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest;                                  // LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> LCD_DMA_Controller_avalon_dma_master_translator:uav_waitrequest
	wire    [1:0] lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount;                                   // LCD_DMA_Controller_avalon_dma_master_translator:uav_burstcount -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata;                                    // LCD_DMA_Controller_avalon_dma_master_translator:uav_writedata -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address;                                      // LCD_DMA_Controller_avalon_dma_master_translator:uav_address -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock;                                         // LCD_DMA_Controller_avalon_dma_master_translator:uav_lock -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write;                                        // LCD_DMA_Controller_avalon_dma_master_translator:uav_write -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read;                                         // LCD_DMA_Controller_avalon_dma_master_translator:uav_read -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata;                                     // LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> LCD_DMA_Controller_avalon_dma_master_translator:uav_readdata
	wire          lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess;                                  // LCD_DMA_Controller_avalon_dma_master_translator:uav_debugaccess -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable;                                   // LCD_DMA_Controller_avalon_dma_master_translator:uav_byteenable -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid;                                // LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> LCD_DMA_Controller_avalon_dma_master_translator:uav_readdatavalid
	wire          vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest;                                  // VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> VGA_DMA_Controller_avalon_dma_master_translator:uav_waitrequest
	wire    [1:0] vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount;                                   // VGA_DMA_Controller_avalon_dma_master_translator:uav_burstcount -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata;                                    // VGA_DMA_Controller_avalon_dma_master_translator:uav_writedata -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address;                                      // VGA_DMA_Controller_avalon_dma_master_translator:uav_address -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock;                                         // VGA_DMA_Controller_avalon_dma_master_translator:uav_lock -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write;                                        // VGA_DMA_Controller_avalon_dma_master_translator:uav_write -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read;                                         // VGA_DMA_Controller_avalon_dma_master_translator:uav_read -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata;                                     // VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> VGA_DMA_Controller_avalon_dma_master_translator:uav_readdata
	wire          vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess;                                  // VGA_DMA_Controller_avalon_dma_master_translator:uav_debugaccess -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable;                                   // VGA_DMA_Controller_avalon_dma_master_translator:uav_byteenable -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid;                                // VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> VGA_DMA_Controller_avalon_dma_master_translator:uav_readdatavalid
	wire          videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_waitrequest;                                 // VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> VideoConferencing_DMA_0_avalon_master_translator:uav_waitrequest
	wire    [1:0] videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_burstcount;                                  // VideoConferencing_DMA_0_avalon_master_translator:uav_burstcount -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_writedata;                                   // VideoConferencing_DMA_0_avalon_master_translator:uav_writedata -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_address;                                     // VideoConferencing_DMA_0_avalon_master_translator:uav_address -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_lock;                                        // VideoConferencing_DMA_0_avalon_master_translator:uav_lock -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_write;                                       // VideoConferencing_DMA_0_avalon_master_translator:uav_write -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_read;                                        // VideoConferencing_DMA_0_avalon_master_translator:uav_read -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_readdata;                                    // VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> VideoConferencing_DMA_0_avalon_master_translator:uav_readdata
	wire          videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_debugaccess;                                 // VideoConferencing_DMA_0_avalon_master_translator:uav_debugaccess -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_byteenable;                                  // VideoConferencing_DMA_0_avalon_master_translator:uav_byteenable -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_readdatavalid;                               // VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> VideoConferencing_DMA_0_avalon_master_translator:uav_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                         // CPU_jtag_debug_module_translator:uav_waitrequest -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                                          // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> CPU_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                                           // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> CPU_jtag_debug_module_translator:uav_writedata
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                             // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> CPU_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                               // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> CPU_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                                // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> CPU_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                                // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> CPU_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                            // CPU_jtag_debug_module_translator:uav_readdata -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                       // CPU_jtag_debug_module_translator:uav_readdatavalid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                         // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CPU_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                                          // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> CPU_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                  // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                                         // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                               // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                     // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                             // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                      // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                     // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                   // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                    // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                   // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                      // SDRAM_s1_translator:uav_waitrequest -> SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                       // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SDRAM_s1_translator:uav_burstcount
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                        // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SDRAM_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                          // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> SDRAM_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                            // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> SDRAM_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                             // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SDRAM_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                             // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> SDRAM_s1_translator:uav_read
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                         // SDRAM_s1_translator:uav_readdata -> SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                    // SDRAM_s1_translator:uav_readdatavalid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                      // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SDRAM_s1_translator:uav_debugaccess
	wire    [3:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                       // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SDRAM_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                               // SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                     // SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                             // SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                      // SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                     // SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                            // SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                  // SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                          // SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                   // SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                  // SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                // SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                 // SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                // SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                              // Flash_flash_data_translator:uav_waitrequest -> Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] flash_flash_data_translator_avalon_universal_slave_0_agent_m0_burstcount;                                               // Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_burstcount -> Flash_flash_data_translator:uav_burstcount
	wire   [31:0] flash_flash_data_translator_avalon_universal_slave_0_agent_m0_writedata;                                                // Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_writedata -> Flash_flash_data_translator:uav_writedata
	wire   [31:0] flash_flash_data_translator_avalon_universal_slave_0_agent_m0_address;                                                  // Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_address -> Flash_flash_data_translator:uav_address
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_m0_write;                                                    // Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_write -> Flash_flash_data_translator:uav_write
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_m0_lock;                                                     // Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_lock -> Flash_flash_data_translator:uav_lock
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_m0_read;                                                     // Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_read -> Flash_flash_data_translator:uav_read
	wire   [31:0] flash_flash_data_translator_avalon_universal_slave_0_agent_m0_readdata;                                                 // Flash_flash_data_translator:uav_readdata -> Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                            // Flash_flash_data_translator:uav_readdatavalid -> Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                              // Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Flash_flash_data_translator:uav_debugaccess
	wire    [3:0] flash_flash_data_translator_avalon_universal_slave_0_agent_m0_byteenable;                                               // Flash_flash_data_translator_avalon_universal_slave_0_agent:m0_byteenable -> Flash_flash_data_translator:uav_byteenable
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                       // Flash_flash_data_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_valid;                                             // Flash_flash_data_translator_avalon_universal_slave_0_agent:rf_source_valid -> Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                     // Flash_flash_data_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_data;                                              // Flash_flash_data_translator_avalon_universal_slave_0_agent:rf_source_data -> Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_ready;                                             // Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Flash_flash_data_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                    // Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Flash_flash_data_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                          // Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Flash_flash_data_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                  // Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Flash_flash_data_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                           // Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Flash_flash_data_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                          // Flash_flash_data_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                        // Flash_flash_data_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Flash_flash_data_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] flash_flash_data_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                         // Flash_flash_data_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Flash_flash_data_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                        // Flash_flash_data_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Flash_flash_data_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // JTAG_UART_avalon_jtag_slave_translator:uav_waitrequest -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> JTAG_UART_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> JTAG_UART_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                                       // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> JTAG_UART_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                                         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> JTAG_UART_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                          // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> JTAG_UART_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                          // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> JTAG_UART_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // JTAG_UART_avalon_jtag_slave_translator:uav_readdata -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // JTAG_UART_avalon_jtag_slave_translator:uav_readdatavalid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> JTAG_UART_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> JTAG_UART_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                             // Interval_Timer_s1_translator:uav_waitrequest -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                              // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Interval_Timer_s1_translator:uav_burstcount
	wire   [31:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                               // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Interval_Timer_s1_translator:uav_writedata
	wire   [31:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                 // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> Interval_Timer_s1_translator:uav_address
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                   // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> Interval_Timer_s1_translator:uav_write
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                    // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Interval_Timer_s1_translator:uav_lock
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                    // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> Interval_Timer_s1_translator:uav_read
	wire   [31:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                // Interval_Timer_s1_translator:uav_readdata -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                           // Interval_Timer_s1_translator:uav_readdatavalid -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                             // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Interval_Timer_s1_translator:uav_debugaccess
	wire    [3:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                              // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Interval_Timer_s1_translator:uav_byteenable
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                      // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                            // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                    // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                             // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                            // Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                   // Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                         // Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                 // Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                          // Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                         // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                       // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                        // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                       // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                           // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                              // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                         // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                       // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                        // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // Red_LEDs_avalon_parallel_port_slave_translator:uav_waitrequest -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Red_LEDs_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                             // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Red_LEDs_avalon_parallel_port_slave_translator:uav_writedata
	wire   [31:0] red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                               // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Red_LEDs_avalon_parallel_port_slave_translator:uav_address
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                                 // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Red_LEDs_avalon_parallel_port_slave_translator:uav_write
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                  // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Red_LEDs_avalon_parallel_port_slave_translator:uav_lock
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                                  // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Red_LEDs_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                              // Red_LEDs_avalon_parallel_port_slave_translator:uav_readdata -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // Red_LEDs_avalon_parallel_port_slave_translator:uav_readdatavalid -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Red_LEDs_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Red_LEDs_avalon_parallel_port_slave_translator:uav_byteenable
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                           // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // Green_LEDs_avalon_parallel_port_slave_translator:uav_waitrequest -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Green_LEDs_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                           // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Green_LEDs_avalon_parallel_port_slave_translator:uav_writedata
	wire   [31:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                             // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Green_LEDs_avalon_parallel_port_slave_translator:uav_address
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                               // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Green_LEDs_avalon_parallel_port_slave_translator:uav_write
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Green_LEDs_avalon_parallel_port_slave_translator:uav_lock
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                                // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Green_LEDs_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                            // Green_LEDs_avalon_parallel_port_slave_translator:uav_readdata -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // Green_LEDs_avalon_parallel_port_slave_translator:uav_readdatavalid -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Green_LEDs_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Green_LEDs_avalon_parallel_port_slave_translator:uav_byteenable
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                         // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // HEX3_HEX0_avalon_parallel_port_slave_translator:uav_waitrequest -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                            // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_writedata
	wire   [31:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                              // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_address
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                                // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_write
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                 // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_lock
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                                 // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                             // HEX3_HEX0_avalon_parallel_port_slave_translator:uav_readdata -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // HEX3_HEX0_avalon_parallel_port_slave_translator:uav_readdatavalid -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> HEX3_HEX0_avalon_parallel_port_slave_translator:uav_byteenable
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                          // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // HEX7_HEX4_avalon_parallel_port_slave_translator:uav_waitrequest -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> HEX7_HEX4_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                            // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> HEX7_HEX4_avalon_parallel_port_slave_translator:uav_writedata
	wire   [31:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                              // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> HEX7_HEX4_avalon_parallel_port_slave_translator:uav_address
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                                // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> HEX7_HEX4_avalon_parallel_port_slave_translator:uav_write
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                 // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> HEX7_HEX4_avalon_parallel_port_slave_translator:uav_lock
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                                 // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> HEX7_HEX4_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                             // HEX7_HEX4_avalon_parallel_port_slave_translator:uav_readdata -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // HEX7_HEX4_avalon_parallel_port_slave_translator:uav_readdatavalid -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> HEX7_HEX4_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> HEX7_HEX4_avalon_parallel_port_slave_translator:uav_byteenable
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                          // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // Slider_Switches_avalon_parallel_port_slave_translator:uav_waitrequest -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Slider_Switches_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                      // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Slider_Switches_avalon_parallel_port_slave_translator:uav_writedata
	wire   [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                        // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Slider_Switches_avalon_parallel_port_slave_translator:uav_address
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                          // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Slider_Switches_avalon_parallel_port_slave_translator:uav_write
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                           // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Slider_Switches_avalon_parallel_port_slave_translator:uav_lock
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                           // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Slider_Switches_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                       // Slider_Switches_avalon_parallel_port_slave_translator:uav_readdata -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // Slider_Switches_avalon_parallel_port_slave_translator:uav_readdatavalid -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Slider_Switches_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Slider_Switches_avalon_parallel_port_slave_translator:uav_byteenable
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                    // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // Pushbuttons_avalon_parallel_port_slave_translator:uav_waitrequest -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Pushbuttons_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Pushbuttons_avalon_parallel_port_slave_translator:uav_writedata
	wire   [31:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Pushbuttons_avalon_parallel_port_slave_translator:uav_address
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Pushbuttons_avalon_parallel_port_slave_translator:uav_write
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Pushbuttons_avalon_parallel_port_slave_translator:uav_lock
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Pushbuttons_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // Pushbuttons_avalon_parallel_port_slave_translator:uav_readdata -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // Pushbuttons_avalon_parallel_port_slave_translator:uav_readdatavalid -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Pushbuttons_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Pushbuttons_avalon_parallel_port_slave_translator:uav_byteenable
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // Expansion_JP5_avalon_parallel_port_slave_translator:uav_waitrequest -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Expansion_JP5_avalon_parallel_port_slave_translator:uav_burstcount
	wire   [31:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Expansion_JP5_avalon_parallel_port_slave_translator:uav_writedata
	wire   [31:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> Expansion_JP5_avalon_parallel_port_slave_translator:uav_address
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> Expansion_JP5_avalon_parallel_port_slave_translator:uav_write
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Expansion_JP5_avalon_parallel_port_slave_translator:uav_lock
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> Expansion_JP5_avalon_parallel_port_slave_translator:uav_read
	wire   [31:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // Expansion_JP5_avalon_parallel_port_slave_translator:uav_readdata -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // Expansion_JP5_avalon_parallel_port_slave_translator:uav_readdatavalid -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Expansion_JP5_avalon_parallel_port_slave_translator:uav_debugaccess
	wire    [3:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Expansion_JP5_avalon_parallel_port_slave_translator:uav_byteenable
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // Serial_Port_avalon_rs232_slave_translator:uav_waitrequest -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Serial_Port_avalon_rs232_slave_translator:uav_burstcount
	wire   [31:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Serial_Port_avalon_rs232_slave_translator:uav_writedata
	wire   [31:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address;                                    // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_address -> Serial_Port_avalon_rs232_slave_translator:uav_address
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write;                                      // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_write -> Serial_Port_avalon_rs232_slave_translator:uav_write
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                       // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Serial_Port_avalon_rs232_slave_translator:uav_lock
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read;                                       // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_read -> Serial_Port_avalon_rs232_slave_translator:uav_read
	wire   [31:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // Serial_Port_avalon_rs232_slave_translator:uav_readdata -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // Serial_Port_avalon_rs232_slave_translator:uav_readdatavalid -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Serial_Port_avalon_rs232_slave_translator:uav_debugaccess
	wire    [3:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Serial_Port_avalon_rs232_slave_translator:uav_byteenable
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // Char_LCD_16x2_avalon_lcd_slave_translator:uav_waitrequest -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Char_LCD_16x2_avalon_lcd_slave_translator:uav_burstcount
	wire    [7:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Char_LCD_16x2_avalon_lcd_slave_translator:uav_writedata
	wire   [31:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address;                                    // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_address -> Char_LCD_16x2_avalon_lcd_slave_translator:uav_address
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write;                                      // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_write -> Char_LCD_16x2_avalon_lcd_slave_translator:uav_write
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                       // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Char_LCD_16x2_avalon_lcd_slave_translator:uav_lock
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read;                                       // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_read -> Char_LCD_16x2_avalon_lcd_slave_translator:uav_read
	wire    [7:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // Char_LCD_16x2_avalon_lcd_slave_translator:uav_readdata -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // Char_LCD_16x2_avalon_lcd_slave_translator:uav_readdatavalid -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Char_LCD_16x2_avalon_lcd_slave_translator:uav_debugaccess
	wire    [0:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Char_LCD_16x2_avalon_lcd_slave_translator:uav_byteenable
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // PS2_Port_avalon_ps2_slave_translator:uav_waitrequest -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> PS2_Port_avalon_ps2_slave_translator:uav_burstcount
	wire   [31:0] ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> PS2_Port_avalon_ps2_slave_translator:uav_writedata
	wire   [31:0] ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address;                                         // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_address -> PS2_Port_avalon_ps2_slave_translator:uav_address
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write;                                           // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_write -> PS2_Port_avalon_ps2_slave_translator:uav_write
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                            // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_lock -> PS2_Port_avalon_ps2_slave_translator:uav_lock
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read;                                            // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_read -> PS2_Port_avalon_ps2_slave_translator:uav_read
	wire   [31:0] ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // PS2_Port_avalon_ps2_slave_translator:uav_readdata -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // PS2_Port_avalon_ps2_slave_translator:uav_readdatavalid -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PS2_Port_avalon_ps2_slave_translator:uav_debugaccess
	wire    [3:0] ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> PS2_Port_avalon_ps2_slave_translator:uav_byteenable
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // SRAM_avalon_sram_slave_translator:uav_waitrequest -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> SRAM_avalon_sram_slave_translator:uav_burstcount
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> SRAM_avalon_sram_slave_translator:uav_writedata
	wire   [31:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                                            // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> SRAM_avalon_sram_slave_translator:uav_address
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                                              // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> SRAM_avalon_sram_slave_translator:uav_write
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                               // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> SRAM_avalon_sram_slave_translator:uav_lock
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                                               // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> SRAM_avalon_sram_slave_translator:uav_read
	wire   [15:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // SRAM_avalon_sram_slave_translator:uav_readdata -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // SRAM_avalon_sram_slave_translator:uav_readdatavalid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SRAM_avalon_sram_slave_translator:uav_debugaccess
	wire    [1:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> SRAM_avalon_sram_slave_translator:uav_byteenable
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [93:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [93:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                  // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                   // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                  // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // VGA_Char_Buffer_avalon_char_control_slave_translator:uav_waitrequest -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_Char_Buffer_avalon_char_control_slave_translator:uav_burstcount
	wire   [31:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_Char_Buffer_avalon_char_control_slave_translator:uav_writedata
	wire   [31:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> VGA_Char_Buffer_avalon_char_control_slave_translator:uav_address
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> VGA_Char_Buffer_avalon_char_control_slave_translator:uav_write
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_Char_Buffer_avalon_char_control_slave_translator:uav_lock
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> VGA_Char_Buffer_avalon_char_control_slave_translator:uav_read
	wire   [31:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // VGA_Char_Buffer_avalon_char_control_slave_translator:uav_readdata -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // VGA_Char_Buffer_avalon_char_control_slave_translator:uav_readdatavalid -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_Char_Buffer_avalon_char_control_slave_translator:uav_debugaccess
	wire    [3:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_Char_Buffer_avalon_char_control_slave_translator:uav_byteenable
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_waitrequest -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_burstcount
	wire    [7:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_writedata
	wire   [31:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_address -> VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_address
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_write -> VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_write
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_lock
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_read -> VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_read
	wire    [7:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_readdata -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_readdatavalid -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_debugaccess
	wire    [0:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_Char_Buffer_avalon_char_buffer_slave_translator:uav_byteenable
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // OnBoard_AV_avalon_av_config_slave_translator:uav_waitrequest -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> OnBoard_AV_avalon_av_config_slave_translator:uav_burstcount
	wire   [31:0] onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                               // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> OnBoard_AV_avalon_av_config_slave_translator:uav_writedata
	wire   [31:0] onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address;                                 // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_address -> OnBoard_AV_avalon_av_config_slave_translator:uav_address
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write;                                   // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_write -> OnBoard_AV_avalon_av_config_slave_translator:uav_write
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                    // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_lock -> OnBoard_AV_avalon_av_config_slave_translator:uav_lock
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read;                                    // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_read -> OnBoard_AV_avalon_av_config_slave_translator:uav_read
	wire   [31:0] onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                // OnBoard_AV_avalon_av_config_slave_translator:uav_readdata -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // OnBoard_AV_avalon_av_config_slave_translator:uav_readdatavalid -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> OnBoard_AV_avalon_av_config_slave_translator:uav_debugaccess
	wire    [3:0] onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> OnBoard_AV_avalon_av_config_slave_translator:uav_byteenable
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                             // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // PS2_Port_Dual_avalon_ps2_slave_translator:uav_waitrequest -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> PS2_Port_Dual_avalon_ps2_slave_translator:uav_burstcount
	wire   [31:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> PS2_Port_Dual_avalon_ps2_slave_translator:uav_writedata
	wire   [31:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address;                                    // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_address -> PS2_Port_Dual_avalon_ps2_slave_translator:uav_address
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write;                                      // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_write -> PS2_Port_Dual_avalon_ps2_slave_translator:uav_write
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                       // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_lock -> PS2_Port_Dual_avalon_ps2_slave_translator:uav_lock
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read;                                       // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_read -> PS2_Port_Dual_avalon_ps2_slave_translator:uav_read
	wire   [31:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // PS2_Port_Dual_avalon_ps2_slave_translator:uav_readdata -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // PS2_Port_Dual_avalon_ps2_slave_translator:uav_readdatavalid -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PS2_Port_Dual_avalon_ps2_slave_translator:uav_debugaccess
	wire    [3:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> PS2_Port_Dual_avalon_ps2_slave_translator:uav_byteenable
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // Audio_avalon_audio_slave_translator:uav_waitrequest -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Audio_avalon_audio_slave_translator:uav_burstcount
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Audio_avalon_audio_slave_translator:uav_writedata
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address;                                          // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_address -> Audio_avalon_audio_slave_translator:uav_address
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write;                                            // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_write -> Audio_avalon_audio_slave_translator:uav_write
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                             // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Audio_avalon_audio_slave_translator:uav_lock
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read;                                             // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_read -> Audio_avalon_audio_slave_translator:uav_read
	wire   [31:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // Audio_avalon_audio_slave_translator:uav_readdata -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // Audio_avalon_audio_slave_translator:uav_readdatavalid -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Audio_avalon_audio_slave_translator:uav_debugaccess
	wire    [3:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Audio_avalon_audio_slave_translator:uav_byteenable
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // Flash_flash_erase_control_translator:uav_waitrequest -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_burstcount -> Flash_flash_erase_control_translator:uav_burstcount
	wire   [31:0] flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_writedata -> Flash_flash_erase_control_translator:uav_writedata
	wire   [31:0] flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_address;                                         // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_address -> Flash_flash_erase_control_translator:uav_address
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_write;                                           // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_write -> Flash_flash_erase_control_translator:uav_write
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_lock;                                            // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_lock -> Flash_flash_erase_control_translator:uav_lock
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_read;                                            // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_read -> Flash_flash_erase_control_translator:uav_read
	wire   [31:0] flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // Flash_flash_erase_control_translator:uav_readdata -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // Flash_flash_erase_control_translator:uav_readdatavalid -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Flash_flash_erase_control_translator:uav_debugaccess
	wire    [3:0] flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:m0_byteenable -> Flash_flash_erase_control_translator:uav_byteenable
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rf_source_valid -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rf_source_data -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // SD_Card_avalon_sdcard_slave_translator:uav_waitrequest -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_Card_avalon_sdcard_slave_translator:uav_burstcount
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_Card_avalon_sdcard_slave_translator:uav_writedata
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address;                                       // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_address -> SD_Card_avalon_sdcard_slave_translator:uav_address
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write;                                         // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_write -> SD_Card_avalon_sdcard_slave_translator:uav_write
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                          // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_lock -> SD_Card_avalon_sdcard_slave_translator:uav_lock
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read;                                          // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_read -> SD_Card_avalon_sdcard_slave_translator:uav_read
	wire   [31:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // SD_Card_avalon_sdcard_slave_translator:uav_readdata -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // SD_Card_avalon_sdcard_slave_translator:uav_readdatavalid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_Card_avalon_sdcard_slave_translator:uav_debugaccess
	wire    [3:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_Card_avalon_sdcard_slave_translator:uav_byteenable
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // IrDA_avalon_irda_slave_translator:uav_waitrequest -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> IrDA_avalon_irda_slave_translator:uav_burstcount
	wire   [31:0] irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> IrDA_avalon_irda_slave_translator:uav_writedata
	wire   [31:0] irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_address;                                            // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_address -> IrDA_avalon_irda_slave_translator:uav_address
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_write;                                              // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_write -> IrDA_avalon_irda_slave_translator:uav_write
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                               // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_lock -> IrDA_avalon_irda_slave_translator:uav_lock
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_read;                                               // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_read -> IrDA_avalon_irda_slave_translator:uav_read
	wire   [31:0] irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // IrDA_avalon_irda_slave_translator:uav_readdata -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // IrDA_avalon_irda_slave_translator:uav_readdatavalid -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> IrDA_avalon_irda_slave_translator:uav_debugaccess
	wire    [3:0] irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> IrDA_avalon_irda_slave_translator:uav_byteenable
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_waitrequest -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_burstcount
	wire   [31:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_writedata
	wire   [31:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_address
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_write
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_lock
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_read
	wire   [31:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_readdata -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_readdatavalid -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_debugaccess
	wire    [3:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Video_In_DMA_Controller_avalon_dma_control_slave_translator:uav_byteenable
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_waitrequest -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_burstcount
	wire   [31:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_writedata
	wire   [31:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_address
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_write
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_lock
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_read
	wire   [31:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_readdata -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_readdatavalid -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_debugaccess
	wire    [3:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Camera_DMA_Controller_avalon_dma_control_slave_translator:uav_byteenable
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // Camera_Config_avalon_av_config_slave_translator:uav_waitrequest -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Camera_Config_avalon_av_config_slave_translator:uav_burstcount
	wire   [31:0] camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                            // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Camera_Config_avalon_av_config_slave_translator:uav_writedata
	wire   [31:0] camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address;                              // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_address -> Camera_Config_avalon_av_config_slave_translator:uav_address
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write;                                // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_write -> Camera_Config_avalon_av_config_slave_translator:uav_write
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                 // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Camera_Config_avalon_av_config_slave_translator:uav_lock
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read;                                 // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_read -> Camera_Config_avalon_av_config_slave_translator:uav_read
	wire   [31:0] camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                             // Camera_Config_avalon_av_config_slave_translator:uav_readdata -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // Camera_Config_avalon_av_config_slave_translator:uav_readdatavalid -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Camera_Config_avalon_av_config_slave_translator:uav_debugaccess
	wire    [3:0] camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Camera_Config_avalon_av_config_slave_translator:uav_byteenable
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                          // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_waitrequest -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_burstcount
	wire    [7:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_writedata
	wire   [31:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_address -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_address
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_write -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_write
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_lock
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_read -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_read
	wire    [7:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_readdata -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_readdatavalid -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_debugaccess
	wire    [0:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator:uav_byteenable
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // USB_avalon_usb_slave_translator:uav_waitrequest -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> USB_avalon_usb_slave_translator:uav_burstcount
	wire   [31:0] usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> USB_avalon_usb_slave_translator:uav_writedata
	wire   [31:0] usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_address;                                              // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_address -> USB_avalon_usb_slave_translator:uav_address
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_write;                                                // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_write -> USB_avalon_usb_slave_translator:uav_write
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_lock -> USB_avalon_usb_slave_translator:uav_lock
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_read;                                                 // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_read -> USB_avalon_usb_slave_translator:uav_read
	wire   [31:0] usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // USB_avalon_usb_slave_translator:uav_readdata -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // USB_avalon_usb_slave_translator:uav_readdatavalid -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> USB_avalon_usb_slave_translator:uav_debugaccess
	wire    [3:0] usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> USB_avalon_usb_slave_translator:uav_byteenable
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // LCD_Char_Buffer_avalon_char_control_slave_translator:uav_waitrequest -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> LCD_Char_Buffer_avalon_char_control_slave_translator:uav_burstcount
	wire   [31:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> LCD_Char_Buffer_avalon_char_control_slave_translator:uav_writedata
	wire   [31:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> LCD_Char_Buffer_avalon_char_control_slave_translator:uav_address
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> LCD_Char_Buffer_avalon_char_control_slave_translator:uav_write
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> LCD_Char_Buffer_avalon_char_control_slave_translator:uav_lock
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> LCD_Char_Buffer_avalon_char_control_slave_translator:uav_read
	wire   [31:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // LCD_Char_Buffer_avalon_char_control_slave_translator:uav_readdata -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // LCD_Char_Buffer_avalon_char_control_slave_translator:uav_readdatavalid -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LCD_Char_Buffer_avalon_char_control_slave_translator:uav_debugaccess
	wire    [3:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> LCD_Char_Buffer_avalon_char_control_slave_translator:uav_byteenable
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_waitrequest -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_burstcount
	wire    [7:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_writedata
	wire   [31:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_address -> LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_address
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_write -> LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_write
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_lock -> LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_lock
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_read -> LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_read
	wire    [7:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_readdata -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_readdatavalid -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_debugaccess
	wire    [0:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> LCD_Char_Buffer_avalon_char_buffer_slave_translator:uav_byteenable
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [84:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [84:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                             // enet_control_port_translator:uav_waitrequest -> enet_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] enet_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                                              // enet_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> enet_control_port_translator:uav_burstcount
	wire   [31:0] enet_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                                               // enet_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> enet_control_port_translator:uav_writedata
	wire   [31:0] enet_control_port_translator_avalon_universal_slave_0_agent_m0_address;                                                 // enet_control_port_translator_avalon_universal_slave_0_agent:m0_address -> enet_control_port_translator:uav_address
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_m0_write;                                                   // enet_control_port_translator_avalon_universal_slave_0_agent:m0_write -> enet_control_port_translator:uav_write
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                                                    // enet_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> enet_control_port_translator:uav_lock
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_m0_read;                                                    // enet_control_port_translator_avalon_universal_slave_0_agent:m0_read -> enet_control_port_translator:uav_read
	wire   [31:0] enet_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                                                // enet_control_port_translator:uav_readdata -> enet_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                           // enet_control_port_translator:uav_readdatavalid -> enet_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                             // enet_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> enet_control_port_translator:uav_debugaccess
	wire    [3:0] enet_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                                              // enet_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> enet_control_port_translator:uav_byteenable
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                      // enet_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;                                            // enet_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                    // enet_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                                             // enet_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;                                            // enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> enet_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                   // enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> enet_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                         // enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> enet_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                 // enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> enet_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                          // enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> enet_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                         // enet_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                       // enet_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> enet_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] enet_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                        // enet_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> enet_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                       // enet_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> enet_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                              // packet_memory_s1_translator:uav_waitrequest -> packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                               // packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> packet_memory_s1_translator:uav_burstcount
	wire   [31:0] packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                // packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> packet_memory_s1_translator:uav_writedata
	wire   [31:0] packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                  // packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> packet_memory_s1_translator:uav_address
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                    // packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> packet_memory_s1_translator:uav_write
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                     // packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> packet_memory_s1_translator:uav_lock
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                     // packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> packet_memory_s1_translator:uav_read
	wire   [31:0] packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                 // packet_memory_s1_translator:uav_readdata -> packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                            // packet_memory_s1_translator:uav_readdatavalid -> packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                              // packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> packet_memory_s1_translator:uav_debugaccess
	wire    [3:0] packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                               // packet_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> packet_memory_s1_translator:uav_byteenable
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                       // packet_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                             // packet_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                     // packet_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                              // packet_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                             // packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> packet_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                    // packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> packet_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                          // packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> packet_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                  // packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> packet_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                           // packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> packet_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                          // packet_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                        // packet_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> packet_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] packet_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                         // packet_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> packet_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                        // packet_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> packet_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // descriptor_memory_s1_translator:uav_waitrequest -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> descriptor_memory_s1_translator:uav_burstcount
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> descriptor_memory_s1_translator:uav_writedata
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                                              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> descriptor_memory_s1_translator:uav_address
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> descriptor_memory_s1_translator:uav_write
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> descriptor_memory_s1_translator:uav_lock
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> descriptor_memory_s1_translator:uav_read
	wire   [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // descriptor_memory_s1_translator:uav_readdata -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // descriptor_memory_s1_translator:uav_readdatavalid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> descriptor_memory_s1_translator:uav_debugaccess
	wire    [3:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> descriptor_memory_s1_translator:uav_byteenable
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_waitrequest -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_burstcount
	wire   [31:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_writedata
	wire   [31:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_address
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_write
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_lock
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_read
	wire   [31:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_readdata -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_readdatavalid -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_debugaccess
	wire    [3:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> LCD_DMA_Controller_avalon_dma_control_slave_translator:uav_byteenable
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_waitrequest -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_burstcount
	wire   [31:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_writedata
	wire   [31:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_address
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_write
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_lock
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_read
	wire   [31:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_readdata -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_readdatavalid -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_debugaccess
	wire    [3:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_DMA_Controller_avalon_dma_control_slave_translator:uav_byteenable
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // VideoConferencing_DMA_0_avalon_slave_translator:uav_waitrequest -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> VideoConferencing_DMA_0_avalon_slave_translator:uav_burstcount
	wire   [31:0] videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                            // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> VideoConferencing_DMA_0_avalon_slave_translator:uav_writedata
	wire   [31:0] videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                              // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> VideoConferencing_DMA_0_avalon_slave_translator:uav_address
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                                // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> VideoConferencing_DMA_0_avalon_slave_translator:uav_write
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                 // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> VideoConferencing_DMA_0_avalon_slave_translator:uav_lock
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                                 // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> VideoConferencing_DMA_0_avalon_slave_translator:uav_read
	wire   [31:0] videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                             // VideoConferencing_DMA_0_avalon_slave_translator:uav_readdata -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // VideoConferencing_DMA_0_avalon_slave_translator:uav_readdatavalid -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VideoConferencing_DMA_0_avalon_slave_translator:uav_debugaccess
	wire    [3:0] videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> VideoConferencing_DMA_0_avalon_slave_translator:uav_byteenable
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [111:0] videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                          // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [111:0] videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                       // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                             // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                     // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [110:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                              // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                             // addr_router:sink_ready -> CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                              // CPU_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                                    // CPU_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                            // CPU_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [110:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                                     // CPU_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                                    // addr_router_001:sink_ready -> CPU_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                    // Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid;                          // Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                  // Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [92:0] video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data;                           // Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready;                          // addr_router_002:sink_ready -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid;                            // Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire   [92:0] camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data;                             // Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_003:sink_ready -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid;                               // LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire   [92:0] lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data;                                // LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router_004:sink_ready -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid;                               // VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire   [92:0] vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data;                                // VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router_005:sink_ready -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	wire          videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                              // VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	wire          videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	wire   [92:0] videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                               // VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	wire          videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_006:sink_ready -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                         // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                               // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                       // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [110:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                                // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                               // id_router:sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                      // SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                            // SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                    // SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [110:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                             // SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                            // id_router_001:sink_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                              // Flash_flash_data_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rp_valid;                                                    // Flash_flash_data_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                            // Flash_flash_data_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [110:0] flash_flash_data_translator_avalon_universal_slave_0_agent_rp_data;                                                     // Flash_flash_data_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          flash_flash_data_translator_avalon_universal_slave_0_agent_rp_ready;                                                    // id_router_002:sink_ready -> Flash_flash_data_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [110:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                          // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_003:sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                             // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                   // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                           // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [110:0] interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                    // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                   // id_router_004:sink_ready -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [110:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                                 // id_router_005:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                 // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [110:0] red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                                  // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_006:sink_ready -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                               // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [110:0] green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                                // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_007:sink_ready -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [110:0] hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                                 // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_008:sink_ready -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [110:0] hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                                 // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_009:sink_ready -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                          // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [110:0] slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                           // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_010:sink_ready -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [110:0] pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_011:sink_ready -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [110:0] expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_012:sink_ready -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                      // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [110:0] serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data;                                       // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_013:sink_ready -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                      // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire   [83:0] char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data;                                       // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_014:sink_ready -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                           // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [110:0] ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data;                                            // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_015:sink_ready -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                              // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire   [92:0] sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                                               // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_016:sink_ready -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [110:0] vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_017:sink_ready -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire   [83:0] vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_018:sink_ready -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                   // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [110:0] onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data;                                    // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_019:sink_ready -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                      // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [110:0] ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data;                                       // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_020:sink_ready -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                            // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [110:0] audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data;                                             // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire          audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_021:sink_ready -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_valid;                                           // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [110:0] flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_data;                                            // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire          flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_022:sink_ready -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                         // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire  [110:0] sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data;                                          // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire          sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_023:sink_ready -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                              // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire  [110:0] irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_data;                                               // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire          irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_024:sink_ready -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire  [110:0] video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire          video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_025:sink_ready -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire  [110:0] camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire          camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_026:sink_ready -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire  [110:0] camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data;                                 // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire          camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_027:sink_ready -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire   [83:0] accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire          accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_028:sink_ready -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                                // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	wire  [110:0] usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_data;                                                 // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	wire          usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_029:sink_ready -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	wire  [110:0] lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	wire          lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_030:sink_ready -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_031:sink_endofpacket
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_031:sink_valid
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_031:sink_startofpacket
	wire   [83:0] lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_031:sink_data
	wire          lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_031:sink_ready -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                             // enet_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_032:sink_endofpacket
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                                                   // enet_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_032:sink_valid
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                           // enet_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_032:sink_startofpacket
	wire  [110:0] enet_control_port_translator_avalon_universal_slave_0_agent_rp_data;                                                    // enet_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_032:sink_data
	wire          enet_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                                                   // id_router_032:sink_ready -> enet_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                              // packet_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_033:sink_endofpacket
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                    // packet_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_033:sink_valid
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                            // packet_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_033:sink_startofpacket
	wire  [110:0] packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                     // packet_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_033:sink_data
	wire          packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                    // id_router_033:sink_ready -> packet_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_034:sink_endofpacket
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_034:sink_valid
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_034:sink_startofpacket
	wire  [110:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_034:sink_data
	wire          descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_034:sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_035:sink_endofpacket
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_035:sink_valid
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_035:sink_startofpacket
	wire  [110:0] lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_035:sink_data
	wire          lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_035:sink_ready -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_036:sink_endofpacket
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_036:sink_valid
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_036:sink_startofpacket
	wire  [110:0] vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_036:sink_data
	wire          vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_036:sink_ready -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_037:sink_endofpacket
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_037:sink_valid
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_037:sink_startofpacket
	wire  [110:0] videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                                 // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_037:sink_data
	wire          videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_037:sink_ready -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                                            // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                                  // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                                          // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [110:0] addr_router_src_data;                                                                                                   // addr_router:src_data -> limiter:cmd_sink_data
	wire   [37:0] addr_router_src_channel;                                                                                                // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                                  // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                                            // limiter:rsp_src_endofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                                  // limiter:rsp_src_valid -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                                          // limiter:rsp_src_startofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [110:0] limiter_rsp_src_data;                                                                                                   // limiter:rsp_src_data -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [37:0] limiter_rsp_src_channel;                                                                                                // limiter:rsp_src_channel -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                                  // CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                                      // burst_adapter:source0_endofpacket -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                            // burst_adapter:source0_valid -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                                    // burst_adapter:source0_startofpacket -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] burst_adapter_source0_data;                                                                                             // burst_adapter:source0_data -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                            // Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [37:0] burst_adapter_source0_channel;                                                                                          // burst_adapter:source0_channel -> Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                                  // burst_adapter_001:source0_endofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                                        // burst_adapter_001:source0_valid -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                                // burst_adapter_001:source0_startofpacket -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [92:0] burst_adapter_001_source0_data;                                                                                         // burst_adapter_001:source0_data -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                                        // SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [37:0] burst_adapter_001_source0_channel;                                                                                      // burst_adapter_001:source0_channel -> SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                                  // burst_adapter_002:source0_endofpacket -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                                        // burst_adapter_002:source0_valid -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                                // burst_adapter_002:source0_startofpacket -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] burst_adapter_002_source0_data;                                                                                         // burst_adapter_002:source0_data -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                                        // VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire   [37:0] burst_adapter_002_source0_channel;                                                                                      // burst_adapter_002:source0_channel -> VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                                                  // burst_adapter_003:source0_endofpacket -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                                        // burst_adapter_003:source0_valid -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                                                // burst_adapter_003:source0_startofpacket -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] burst_adapter_003_source0_data;                                                                                         // burst_adapter_003:source0_data -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                                        // Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire   [37:0] burst_adapter_003_source0_channel;                                                                                      // burst_adapter_003:source0_channel -> Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_004_source0_endofpacket;                                                                                  // burst_adapter_004:source0_endofpacket -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_004_source0_valid;                                                                                        // burst_adapter_004:source0_valid -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_004_source0_startofpacket;                                                                                // burst_adapter_004:source0_startofpacket -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [83:0] burst_adapter_004_source0_data;                                                                                         // burst_adapter_004:source0_data -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_004_source0_ready;                                                                                        // LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_004:source0_ready
	wire   [37:0] burst_adapter_004_source0_channel;                                                                                      // burst_adapter_004:source0_channel -> LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                         // rst_controller:reset_out -> [Accelerometer:reset, Accelerometer_avalon_accelerometer_spi_mode_slave_translator:reset, Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent:reset, Accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Audio:reset, Audio_avalon_audio_slave_translator:reset, Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:reset, Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CPU:reset_n, CPU_data_master_translator:reset, CPU_data_master_translator_avalon_universal_master_0_agent:reset, CPU_instruction_master_translator:reset, CPU_instruction_master_translator_avalon_universal_master_0_agent:reset, CPU_jtag_debug_module_translator:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Camera_Bayer_Resampler:reset, Camera_Clipper:reset, Camera_Config:reset, Camera_Config_avalon_av_config_slave_translator:reset, Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:reset, Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Camera_DMA_Controller:reset, Camera_DMA_Controller_avalon_dma_control_slave_translator:reset, Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:reset, Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Camera_DMA_Controller_avalon_dma_master_translator:reset, Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:reset, Camera_In:reset, Camera_RGB_Resampler:reset, Camera_Scaler:reset, Char_LCD_16x2:reset, Char_LCD_16x2_avalon_lcd_slave_translator:reset, Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:reset, Char_LCD_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Expansion_JP5:reset, Expansion_JP5_avalon_parallel_port_slave_translator:reset, Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Green_LEDs:reset, Green_LEDs_avalon_parallel_port_slave_translator:reset, Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, HEX3_HEX0:reset, HEX3_HEX0_avalon_parallel_port_slave_translator:reset, HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, HEX7_HEX4:reset, HEX7_HEX4_avalon_parallel_port_slave_translator:reset, HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Interval_Timer:reset_n, Interval_Timer_s1_translator:reset, Interval_Timer_s1_translator_avalon_universal_slave_0_agent:reset, Interval_Timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, JTAG_UART:rst_n, JTAG_UART_avalon_jtag_slave_translator:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LCD_Alpha_Blender:reset, LCD_Char_Buffer:reset, LCD_Char_Buffer_avalon_char_buffer_slave_translator:reset, LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:reset, LCD_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LCD_Char_Buffer_avalon_char_control_slave_translator:reset, LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:reset, LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LCD_Dual_Clock_FIFO:reset_stream_in, LCD_RGB_Resampler:reset, LCD_Scalar:reset, OnBoard_AV:reset, OnBoard_AV_avalon_av_config_slave_translator:reset, OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:reset, OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, PS2_Port:reset, PS2_Port_Dual:reset, PS2_Port_Dual_avalon_ps2_slave_translator:reset, PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:reset, PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, PS2_Port_avalon_ps2_slave_translator:reset, PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:reset, PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Pushbuttons:reset, Pushbuttons_avalon_parallel_port_slave_translator:reset, Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Red_LEDs:reset, Red_LEDs_avalon_parallel_port_slave_translator:reset, Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SDRAM:reset_n, SDRAM_s1_translator:reset, SDRAM_s1_translator_avalon_universal_slave_0_agent:reset, SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SRAM:reset, SRAM_avalon_sram_slave_translator:reset, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, SRAM_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Serial_Port:reset, Serial_Port_avalon_rs232_slave_translator:reset, Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:reset, Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Slider_Switches:reset, Slider_Switches_avalon_parallel_port_slave_translator:reset, Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, USB:reset, USB_avalon_usb_slave_translator:reset, USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:reset, USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Alpha_Blender:reset, VGA_Char_Buffer:reset, VGA_Char_Buffer_avalon_char_buffer_slave_translator:reset, VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:reset, VGA_Char_Buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Char_Buffer_avalon_char_control_slave_translator:reset, VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:reset, VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_Dual_Clock_FIFO:reset_stream_in, VGA_Pixel_RGB_Resampler:reset, VGA_Pixel_Scaler:reset, Video_In:reset, Video_In_CSC:reset, Video_In_Chroma_Resampler:reset, Video_In_Clipper:reset, Video_In_DMA_Controller:reset, Video_In_DMA_Controller_avalon_dma_control_slave_translator:reset, Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:reset, Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Video_In_DMA_Controller_avalon_dma_master_translator:reset, Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:reset, Video_In_RGB_Resampler:reset, Video_In_Scaler:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, burst_adapter_004:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_016:reset, id_router:reset, id_router_001:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_025:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, id_router_029:reset, id_router_030:reset, id_router_031:reset, irq_mapper:reset, limiter:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_demux_029:reset, rsp_xbar_demux_030:reset, rsp_xbar_demux_031:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset]
	wire          rst_controller_001_reset_out_reset;                                                                                     // rst_controller_001:reset_out -> [VGA_Controller:reset, VGA_Dual_Clock_FIFO:reset_stream_out]
	wire          rst_controller_002_reset_out_reset;                                                                                     // rst_controller_002:reset_out -> External_Clocks:reset
	wire          rst_controller_003_reset_out_reset;                                                                                     // rst_controller_003:reset_out -> [Flash:i_reset_n, Flash_flash_data_translator:reset, Flash_flash_data_translator_avalon_universal_slave_0_agent:reset, Flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Flash_flash_erase_control_translator:reset, Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:reset, Flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, IrDA:reset, IrDA_avalon_irda_slave_translator:reset, IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:reset, IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_Card:i_reset_n, SD_Card_avalon_sdcard_slave_translator:reset, SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:reset, SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_002:reset, id_router_002:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset]
	wire          rst_controller_004_reset_out_reset;                                                                                     // rst_controller_004:reset_out -> [LCD_Controller:reset, LCD_Dual_Clock_FIFO:reset_stream_out]
	wire          rst_controller_005_reset_out_reset;                                                                                     // rst_controller_005:reset_out -> [avalon_st_adapter:in_rst_0_reset, descriptor_memory:reset, descriptor_memory_s1_translator:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, enet:reset, enet_control_port_translator:reset, enet_control_port_translator_avalon_universal_slave_0_agent:reset, enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_032:reset, id_router_033:reset, id_router_034:reset, packet_memory:reset, packet_memory_s1_translator:reset, packet_memory_s1_translator_avalon_universal_slave_0_agent:reset, packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_032:reset, rsp_xbar_demux_033:reset, rsp_xbar_demux_034:reset]
	wire          rst_controller_005_reset_out_reset_req;                                                                                 // rst_controller_005:reset_req -> [descriptor_memory:reset_req, packet_memory:reset_req]
	wire          rst_controller_006_reset_out_reset;                                                                                     // rst_controller_006:reset_out -> [VideoConferencing_DMA_0:resetn, VideoConferencing_DMA_0_avalon_master_translator:reset, VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:reset, VideoConferencing_DMA_0_avalon_slave_translator:reset, VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:reset, VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router_006:reset, avalon_st_adapter_001:in_rst_0_reset, cmd_xbar_demux_006:reset, id_router_037:reset, rsp_xbar_demux_037:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                        // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                              // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                                      // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [110:0] cmd_xbar_demux_src0_data;                                                                                               // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [37:0] cmd_xbar_demux_src0_channel;                                                                                            // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                              // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                        // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                              // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                                      // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [110:0] cmd_xbar_demux_src1_data;                                                                                               // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [37:0] cmd_xbar_demux_src1_channel;                                                                                            // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                              // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                                        // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                              // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                                      // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [110:0] cmd_xbar_demux_src2_data;                                                                                               // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [37:0] cmd_xbar_demux_src2_channel;                                                                                            // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                              // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                                    // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                          // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                                  // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src0_data;                                                                                           // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [37:0] cmd_xbar_demux_001_src0_channel;                                                                                        // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                          // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                                    // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                          // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                                  // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src1_data;                                                                                           // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [37:0] cmd_xbar_demux_001_src1_channel;                                                                                        // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                          // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                                    // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                          // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                                  // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src2_data;                                                                                           // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [37:0] cmd_xbar_demux_001_src2_channel;                                                                                        // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                                          // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                                    // cmd_xbar_demux_001:src3_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                          // cmd_xbar_demux_001:src3_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                                  // cmd_xbar_demux_001:src3_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src3_data;                                                                                           // cmd_xbar_demux_001:src3_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src3_channel;                                                                                        // cmd_xbar_demux_001:src3_channel -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                                    // cmd_xbar_demux_001:src4_endofpacket -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                          // cmd_xbar_demux_001:src4_valid -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                                  // cmd_xbar_demux_001:src4_startofpacket -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src4_data;                                                                                           // cmd_xbar_demux_001:src4_data -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src4_channel;                                                                                        // cmd_xbar_demux_001:src4_channel -> Interval_Timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                                    // cmd_xbar_demux_001:src5_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                                          // cmd_xbar_demux_001:src5_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                                  // cmd_xbar_demux_001:src5_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src5_data;                                                                                           // cmd_xbar_demux_001:src5_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src5_channel;                                                                                        // cmd_xbar_demux_001:src5_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                                    // cmd_xbar_demux_001:src6_endofpacket -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                                          // cmd_xbar_demux_001:src6_valid -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                                  // cmd_xbar_demux_001:src6_startofpacket -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src6_data;                                                                                           // cmd_xbar_demux_001:src6_data -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src6_channel;                                                                                        // cmd_xbar_demux_001:src6_channel -> Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                                    // cmd_xbar_demux_001:src7_endofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                                          // cmd_xbar_demux_001:src7_valid -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                                  // cmd_xbar_demux_001:src7_startofpacket -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src7_data;                                                                                           // cmd_xbar_demux_001:src7_data -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src7_channel;                                                                                        // cmd_xbar_demux_001:src7_channel -> Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                                    // cmd_xbar_demux_001:src8_endofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                                          // cmd_xbar_demux_001:src8_valid -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                                  // cmd_xbar_demux_001:src8_startofpacket -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src8_data;                                                                                           // cmd_xbar_demux_001:src8_data -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src8_channel;                                                                                        // cmd_xbar_demux_001:src8_channel -> HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                                    // cmd_xbar_demux_001:src9_endofpacket -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                                          // cmd_xbar_demux_001:src9_valid -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                                  // cmd_xbar_demux_001:src9_startofpacket -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src9_data;                                                                                           // cmd_xbar_demux_001:src9_data -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src9_channel;                                                                                        // cmd_xbar_demux_001:src9_channel -> HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                                   // cmd_xbar_demux_001:src10_endofpacket -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                                         // cmd_xbar_demux_001:src10_valid -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                                 // cmd_xbar_demux_001:src10_startofpacket -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src10_data;                                                                                          // cmd_xbar_demux_001:src10_data -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src10_channel;                                                                                       // cmd_xbar_demux_001:src10_channel -> Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                                   // cmd_xbar_demux_001:src11_endofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                                         // cmd_xbar_demux_001:src11_valid -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                                 // cmd_xbar_demux_001:src11_startofpacket -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src11_data;                                                                                          // cmd_xbar_demux_001:src11_data -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src11_channel;                                                                                       // cmd_xbar_demux_001:src11_channel -> Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                                   // cmd_xbar_demux_001:src12_endofpacket -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                                         // cmd_xbar_demux_001:src12_valid -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                                 // cmd_xbar_demux_001:src12_startofpacket -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src12_data;                                                                                          // cmd_xbar_demux_001:src12_data -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src12_channel;                                                                                       // cmd_xbar_demux_001:src12_channel -> Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                                                   // cmd_xbar_demux_001:src13_endofpacket -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                                         // cmd_xbar_demux_001:src13_valid -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                                                 // cmd_xbar_demux_001:src13_startofpacket -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src13_data;                                                                                          // cmd_xbar_demux_001:src13_data -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src13_channel;                                                                                       // cmd_xbar_demux_001:src13_channel -> Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                                                   // cmd_xbar_demux_001:src15_endofpacket -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                                         // cmd_xbar_demux_001:src15_valid -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                                                 // cmd_xbar_demux_001:src15_startofpacket -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src15_data;                                                                                          // cmd_xbar_demux_001:src15_data -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src15_channel;                                                                                       // cmd_xbar_demux_001:src15_channel -> PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src17_endofpacket;                                                                                   // cmd_xbar_demux_001:src17_endofpacket -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src17_valid;                                                                                         // cmd_xbar_demux_001:src17_valid -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src17_startofpacket;                                                                                 // cmd_xbar_demux_001:src17_startofpacket -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src17_data;                                                                                          // cmd_xbar_demux_001:src17_data -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src17_channel;                                                                                       // cmd_xbar_demux_001:src17_channel -> VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src19_endofpacket;                                                                                   // cmd_xbar_demux_001:src19_endofpacket -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src19_valid;                                                                                         // cmd_xbar_demux_001:src19_valid -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src19_startofpacket;                                                                                 // cmd_xbar_demux_001:src19_startofpacket -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src19_data;                                                                                          // cmd_xbar_demux_001:src19_data -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src19_channel;                                                                                       // cmd_xbar_demux_001:src19_channel -> OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src20_endofpacket;                                                                                   // cmd_xbar_demux_001:src20_endofpacket -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src20_valid;                                                                                         // cmd_xbar_demux_001:src20_valid -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src20_startofpacket;                                                                                 // cmd_xbar_demux_001:src20_startofpacket -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src20_data;                                                                                          // cmd_xbar_demux_001:src20_data -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src20_channel;                                                                                       // cmd_xbar_demux_001:src20_channel -> PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src21_endofpacket;                                                                                   // cmd_xbar_demux_001:src21_endofpacket -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src21_valid;                                                                                         // cmd_xbar_demux_001:src21_valid -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src21_startofpacket;                                                                                 // cmd_xbar_demux_001:src21_startofpacket -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src21_data;                                                                                          // cmd_xbar_demux_001:src21_data -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src21_channel;                                                                                       // cmd_xbar_demux_001:src21_channel -> Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src22_endofpacket;                                                                                   // cmd_xbar_demux_001:src22_endofpacket -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src22_valid;                                                                                         // cmd_xbar_demux_001:src22_valid -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src22_startofpacket;                                                                                 // cmd_xbar_demux_001:src22_startofpacket -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src22_data;                                                                                          // cmd_xbar_demux_001:src22_data -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src22_channel;                                                                                       // cmd_xbar_demux_001:src22_channel -> Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src23_endofpacket;                                                                                   // cmd_xbar_demux_001:src23_endofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src23_valid;                                                                                         // cmd_xbar_demux_001:src23_valid -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src23_startofpacket;                                                                                 // cmd_xbar_demux_001:src23_startofpacket -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src23_data;                                                                                          // cmd_xbar_demux_001:src23_data -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src23_channel;                                                                                       // cmd_xbar_demux_001:src23_channel -> SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src24_endofpacket;                                                                                   // cmd_xbar_demux_001:src24_endofpacket -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src24_valid;                                                                                         // cmd_xbar_demux_001:src24_valid -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src24_startofpacket;                                                                                 // cmd_xbar_demux_001:src24_startofpacket -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src24_data;                                                                                          // cmd_xbar_demux_001:src24_data -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src24_channel;                                                                                       // cmd_xbar_demux_001:src24_channel -> IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src25_endofpacket;                                                                                   // cmd_xbar_demux_001:src25_endofpacket -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src25_valid;                                                                                         // cmd_xbar_demux_001:src25_valid -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src25_startofpacket;                                                                                 // cmd_xbar_demux_001:src25_startofpacket -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src25_data;                                                                                          // cmd_xbar_demux_001:src25_data -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src25_channel;                                                                                       // cmd_xbar_demux_001:src25_channel -> Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src26_endofpacket;                                                                                   // cmd_xbar_demux_001:src26_endofpacket -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src26_valid;                                                                                         // cmd_xbar_demux_001:src26_valid -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src26_startofpacket;                                                                                 // cmd_xbar_demux_001:src26_startofpacket -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src26_data;                                                                                          // cmd_xbar_demux_001:src26_data -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src26_channel;                                                                                       // cmd_xbar_demux_001:src26_channel -> Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src27_endofpacket;                                                                                   // cmd_xbar_demux_001:src27_endofpacket -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src27_valid;                                                                                         // cmd_xbar_demux_001:src27_valid -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src27_startofpacket;                                                                                 // cmd_xbar_demux_001:src27_startofpacket -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src27_data;                                                                                          // cmd_xbar_demux_001:src27_data -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src27_channel;                                                                                       // cmd_xbar_demux_001:src27_channel -> Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src29_endofpacket;                                                                                   // cmd_xbar_demux_001:src29_endofpacket -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src29_valid;                                                                                         // cmd_xbar_demux_001:src29_valid -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src29_startofpacket;                                                                                 // cmd_xbar_demux_001:src29_startofpacket -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src29_data;                                                                                          // cmd_xbar_demux_001:src29_data -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src29_channel;                                                                                       // cmd_xbar_demux_001:src29_channel -> USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src30_endofpacket;                                                                                   // cmd_xbar_demux_001:src30_endofpacket -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src30_valid;                                                                                         // cmd_xbar_demux_001:src30_valid -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src30_startofpacket;                                                                                 // cmd_xbar_demux_001:src30_startofpacket -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src30_data;                                                                                          // cmd_xbar_demux_001:src30_data -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src30_channel;                                                                                       // cmd_xbar_demux_001:src30_channel -> LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src32_endofpacket;                                                                                   // cmd_xbar_demux_001:src32_endofpacket -> enet_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src32_valid;                                                                                         // cmd_xbar_demux_001:src32_valid -> enet_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src32_startofpacket;                                                                                 // cmd_xbar_demux_001:src32_startofpacket -> enet_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src32_data;                                                                                          // cmd_xbar_demux_001:src32_data -> enet_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src32_channel;                                                                                       // cmd_xbar_demux_001:src32_channel -> enet_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src33_endofpacket;                                                                                   // cmd_xbar_demux_001:src33_endofpacket -> packet_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src33_valid;                                                                                         // cmd_xbar_demux_001:src33_valid -> packet_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src33_startofpacket;                                                                                 // cmd_xbar_demux_001:src33_startofpacket -> packet_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src33_data;                                                                                          // cmd_xbar_demux_001:src33_data -> packet_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src33_channel;                                                                                       // cmd_xbar_demux_001:src33_channel -> packet_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src34_endofpacket;                                                                                   // cmd_xbar_demux_001:src34_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src34_valid;                                                                                         // cmd_xbar_demux_001:src34_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src34_startofpacket;                                                                                 // cmd_xbar_demux_001:src34_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src34_data;                                                                                          // cmd_xbar_demux_001:src34_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src34_channel;                                                                                       // cmd_xbar_demux_001:src34_channel -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src35_endofpacket;                                                                                   // cmd_xbar_demux_001:src35_endofpacket -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src35_valid;                                                                                         // cmd_xbar_demux_001:src35_valid -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src35_startofpacket;                                                                                 // cmd_xbar_demux_001:src35_startofpacket -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src35_data;                                                                                          // cmd_xbar_demux_001:src35_data -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src35_channel;                                                                                       // cmd_xbar_demux_001:src35_channel -> LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src36_endofpacket;                                                                                   // cmd_xbar_demux_001:src36_endofpacket -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src36_valid;                                                                                         // cmd_xbar_demux_001:src36_valid -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src36_startofpacket;                                                                                 // cmd_xbar_demux_001:src36_startofpacket -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src36_data;                                                                                          // cmd_xbar_demux_001:src36_data -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src36_channel;                                                                                       // cmd_xbar_demux_001:src36_channel -> VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src37_endofpacket;                                                                                   // cmd_xbar_demux_001:src37_endofpacket -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src37_valid;                                                                                         // cmd_xbar_demux_001:src37_valid -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src37_startofpacket;                                                                                 // cmd_xbar_demux_001:src37_startofpacket -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src37_data;                                                                                          // cmd_xbar_demux_001:src37_data -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_demux_001_src37_channel;                                                                                       // cmd_xbar_demux_001:src37_channel -> VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                                    // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_016:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                                          // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_016:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                                  // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_016:sink1_startofpacket
	wire   [92:0] cmd_xbar_demux_002_src0_data;                                                                                           // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_016:sink1_data
	wire   [37:0] cmd_xbar_demux_002_src0_channel;                                                                                        // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_016:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                                          // cmd_xbar_mux_016:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                                    // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_016:sink2_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                                          // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_016:sink2_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                                  // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_016:sink2_startofpacket
	wire   [92:0] cmd_xbar_demux_003_src0_data;                                                                                           // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_016:sink2_data
	wire   [37:0] cmd_xbar_demux_003_src0_channel;                                                                                        // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_016:sink2_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                                          // cmd_xbar_mux_016:sink2_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                                    // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_016:sink3_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                                          // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_016:sink3_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                                                  // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_016:sink3_startofpacket
	wire   [92:0] cmd_xbar_demux_004_src0_data;                                                                                           // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_016:sink3_data
	wire   [37:0] cmd_xbar_demux_004_src0_channel;                                                                                        // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_016:sink3_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                                          // cmd_xbar_mux_016:sink3_ready -> cmd_xbar_demux_004:src0_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                                    // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_016:sink4_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                                          // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_016:sink4_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                                                  // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_016:sink4_startofpacket
	wire   [92:0] cmd_xbar_demux_005_src0_data;                                                                                           // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_016:sink4_data
	wire   [37:0] cmd_xbar_demux_005_src0_channel;                                                                                        // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_016:sink4_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                                          // cmd_xbar_mux_016:sink4_ready -> cmd_xbar_demux_005:src0_ready
	wire          cmd_xbar_demux_006_src0_endofpacket;                                                                                    // cmd_xbar_demux_006:src0_endofpacket -> cmd_xbar_mux_016:sink5_endofpacket
	wire          cmd_xbar_demux_006_src0_valid;                                                                                          // cmd_xbar_demux_006:src0_valid -> cmd_xbar_mux_016:sink5_valid
	wire          cmd_xbar_demux_006_src0_startofpacket;                                                                                  // cmd_xbar_demux_006:src0_startofpacket -> cmd_xbar_mux_016:sink5_startofpacket
	wire   [92:0] cmd_xbar_demux_006_src0_data;                                                                                           // cmd_xbar_demux_006:src0_data -> cmd_xbar_mux_016:sink5_data
	wire   [37:0] cmd_xbar_demux_006_src0_channel;                                                                                        // cmd_xbar_demux_006:src0_channel -> cmd_xbar_mux_016:sink5_channel
	wire          cmd_xbar_demux_006_src0_ready;                                                                                          // cmd_xbar_mux_016:sink5_ready -> cmd_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                        // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                              // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                                      // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [110:0] rsp_xbar_demux_src0_data;                                                                                               // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [37:0] rsp_xbar_demux_src0_channel;                                                                                            // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                              // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                        // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                              // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                                      // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [110:0] rsp_xbar_demux_src1_data;                                                                                               // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [37:0] rsp_xbar_demux_src1_channel;                                                                                            // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                              // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                                    // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                          // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                                  // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [110:0] rsp_xbar_demux_001_src0_data;                                                                                           // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [37:0] rsp_xbar_demux_001_src0_channel;                                                                                        // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                          // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                                    // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                          // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                                  // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [110:0] rsp_xbar_demux_001_src1_data;                                                                                           // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [37:0] rsp_xbar_demux_001_src1_channel;                                                                                        // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                                          // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                                    // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                          // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                                  // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [110:0] rsp_xbar_demux_002_src0_data;                                                                                           // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [37:0] rsp_xbar_demux_002_src0_channel;                                                                                        // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                          // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                                    // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                                          // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                                  // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [110:0] rsp_xbar_demux_002_src1_data;                                                                                           // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [37:0] rsp_xbar_demux_002_src1_channel;                                                                                        // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                                          // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                                    // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                          // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                                  // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [110:0] rsp_xbar_demux_003_src0_data;                                                                                           // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [37:0] rsp_xbar_demux_003_src0_channel;                                                                                        // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                          // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                                    // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                          // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                                  // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [110:0] rsp_xbar_demux_004_src0_data;                                                                                           // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [37:0] rsp_xbar_demux_004_src0_channel;                                                                                        // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                          // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                                    // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                          // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                                  // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [110:0] rsp_xbar_demux_005_src0_data;                                                                                           // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [37:0] rsp_xbar_demux_005_src0_channel;                                                                                        // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                          // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                                    // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                          // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                                  // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [110:0] rsp_xbar_demux_006_src0_data;                                                                                           // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [37:0] rsp_xbar_demux_006_src0_channel;                                                                                        // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                          // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                                    // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                          // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                                  // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [110:0] rsp_xbar_demux_007_src0_data;                                                                                           // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [37:0] rsp_xbar_demux_007_src0_channel;                                                                                        // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                          // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                                    // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                          // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                                  // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [110:0] rsp_xbar_demux_008_src0_data;                                                                                           // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [37:0] rsp_xbar_demux_008_src0_channel;                                                                                        // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                          // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                                    // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                          // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                                  // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [110:0] rsp_xbar_demux_009_src0_data;                                                                                           // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [37:0] rsp_xbar_demux_009_src0_channel;                                                                                        // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                          // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                                    // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                          // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                                  // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [110:0] rsp_xbar_demux_010_src0_data;                                                                                           // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [37:0] rsp_xbar_demux_010_src0_channel;                                                                                        // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                          // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                                    // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                          // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                                  // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [110:0] rsp_xbar_demux_011_src0_data;                                                                                           // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [37:0] rsp_xbar_demux_011_src0_channel;                                                                                        // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                          // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                                    // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                          // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                                  // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [110:0] rsp_xbar_demux_012_src0_data;                                                                                           // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [37:0] rsp_xbar_demux_012_src0_channel;                                                                                        // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                                          // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                                    // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                          // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                                  // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [110:0] rsp_xbar_demux_013_src0_data;                                                                                           // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire   [37:0] rsp_xbar_demux_013_src0_channel;                                                                                        // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                                          // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                                    // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                                          // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                                  // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [110:0] rsp_xbar_demux_015_src0_data;                                                                                           // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire   [37:0] rsp_xbar_demux_015_src0_channel;                                                                                        // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                                          // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src1_endofpacket;                                                                                    // rsp_xbar_demux_016:src1_endofpacket -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_016_src1_valid;                                                                                          // rsp_xbar_demux_016:src1_valid -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_016_src1_startofpacket;                                                                                  // rsp_xbar_demux_016:src1_startofpacket -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [92:0] rsp_xbar_demux_016_src1_data;                                                                                           // rsp_xbar_demux_016:src1_data -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [37:0] rsp_xbar_demux_016_src1_channel;                                                                                        // rsp_xbar_demux_016:src1_channel -> Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_016_src2_endofpacket;                                                                                    // rsp_xbar_demux_016:src2_endofpacket -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_016_src2_valid;                                                                                          // rsp_xbar_demux_016:src2_valid -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_016_src2_startofpacket;                                                                                  // rsp_xbar_demux_016:src2_startofpacket -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [92:0] rsp_xbar_demux_016_src2_data;                                                                                           // rsp_xbar_demux_016:src2_data -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [37:0] rsp_xbar_demux_016_src2_channel;                                                                                        // rsp_xbar_demux_016:src2_channel -> Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_016_src3_endofpacket;                                                                                    // rsp_xbar_demux_016:src3_endofpacket -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_016_src3_valid;                                                                                          // rsp_xbar_demux_016:src3_valid -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_016_src3_startofpacket;                                                                                  // rsp_xbar_demux_016:src3_startofpacket -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [92:0] rsp_xbar_demux_016_src3_data;                                                                                           // rsp_xbar_demux_016:src3_data -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [37:0] rsp_xbar_demux_016_src3_channel;                                                                                        // rsp_xbar_demux_016:src3_channel -> LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_016_src4_endofpacket;                                                                                    // rsp_xbar_demux_016:src4_endofpacket -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_016_src4_valid;                                                                                          // rsp_xbar_demux_016:src4_valid -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_016_src4_startofpacket;                                                                                  // rsp_xbar_demux_016:src4_startofpacket -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [92:0] rsp_xbar_demux_016_src4_data;                                                                                           // rsp_xbar_demux_016:src4_data -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [37:0] rsp_xbar_demux_016_src4_channel;                                                                                        // rsp_xbar_demux_016:src4_channel -> VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_016_src5_endofpacket;                                                                                    // rsp_xbar_demux_016:src5_endofpacket -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_016_src5_valid;                                                                                          // rsp_xbar_demux_016:src5_valid -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_016_src5_startofpacket;                                                                                  // rsp_xbar_demux_016:src5_startofpacket -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [92:0] rsp_xbar_demux_016_src5_data;                                                                                           // rsp_xbar_demux_016:src5_data -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [37:0] rsp_xbar_demux_016_src5_channel;                                                                                        // rsp_xbar_demux_016:src5_channel -> VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                                    // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                                          // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                                  // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [110:0] rsp_xbar_demux_017_src0_data;                                                                                           // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire   [37:0] rsp_xbar_demux_017_src0_channel;                                                                                        // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                                          // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                                                    // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                                          // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                                                  // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [110:0] rsp_xbar_demux_019_src0_data;                                                                                           // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	wire   [37:0] rsp_xbar_demux_019_src0_channel;                                                                                        // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                                          // rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                                                    // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                                          // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                                                  // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	wire  [110:0] rsp_xbar_demux_020_src0_data;                                                                                           // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	wire   [37:0] rsp_xbar_demux_020_src0_channel;                                                                                        // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                                          // rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire          rsp_xbar_demux_021_src0_endofpacket;                                                                                    // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	wire          rsp_xbar_demux_021_src0_valid;                                                                                          // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	wire          rsp_xbar_demux_021_src0_startofpacket;                                                                                  // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	wire  [110:0] rsp_xbar_demux_021_src0_data;                                                                                           // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	wire   [37:0] rsp_xbar_demux_021_src0_channel;                                                                                        // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	wire          rsp_xbar_demux_021_src0_ready;                                                                                          // rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	wire          rsp_xbar_demux_022_src0_endofpacket;                                                                                    // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	wire          rsp_xbar_demux_022_src0_valid;                                                                                          // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink22_valid
	wire          rsp_xbar_demux_022_src0_startofpacket;                                                                                  // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	wire  [110:0] rsp_xbar_demux_022_src0_data;                                                                                           // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink22_data
	wire   [37:0] rsp_xbar_demux_022_src0_channel;                                                                                        // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink22_channel
	wire          rsp_xbar_demux_022_src0_ready;                                                                                          // rsp_xbar_mux_001:sink22_ready -> rsp_xbar_demux_022:src0_ready
	wire          rsp_xbar_demux_023_src0_endofpacket;                                                                                    // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_001:sink23_endofpacket
	wire          rsp_xbar_demux_023_src0_valid;                                                                                          // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_001:sink23_valid
	wire          rsp_xbar_demux_023_src0_startofpacket;                                                                                  // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_001:sink23_startofpacket
	wire  [110:0] rsp_xbar_demux_023_src0_data;                                                                                           // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_001:sink23_data
	wire   [37:0] rsp_xbar_demux_023_src0_channel;                                                                                        // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_001:sink23_channel
	wire          rsp_xbar_demux_023_src0_ready;                                                                                          // rsp_xbar_mux_001:sink23_ready -> rsp_xbar_demux_023:src0_ready
	wire          rsp_xbar_demux_024_src0_endofpacket;                                                                                    // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_001:sink24_endofpacket
	wire          rsp_xbar_demux_024_src0_valid;                                                                                          // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_001:sink24_valid
	wire          rsp_xbar_demux_024_src0_startofpacket;                                                                                  // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_001:sink24_startofpacket
	wire  [110:0] rsp_xbar_demux_024_src0_data;                                                                                           // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_001:sink24_data
	wire   [37:0] rsp_xbar_demux_024_src0_channel;                                                                                        // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_001:sink24_channel
	wire          rsp_xbar_demux_024_src0_ready;                                                                                          // rsp_xbar_mux_001:sink24_ready -> rsp_xbar_demux_024:src0_ready
	wire          rsp_xbar_demux_025_src0_endofpacket;                                                                                    // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_001:sink25_endofpacket
	wire          rsp_xbar_demux_025_src0_valid;                                                                                          // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_001:sink25_valid
	wire          rsp_xbar_demux_025_src0_startofpacket;                                                                                  // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_001:sink25_startofpacket
	wire  [110:0] rsp_xbar_demux_025_src0_data;                                                                                           // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_001:sink25_data
	wire   [37:0] rsp_xbar_demux_025_src0_channel;                                                                                        // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_001:sink25_channel
	wire          rsp_xbar_demux_025_src0_ready;                                                                                          // rsp_xbar_mux_001:sink25_ready -> rsp_xbar_demux_025:src0_ready
	wire          rsp_xbar_demux_026_src0_endofpacket;                                                                                    // rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_001:sink26_endofpacket
	wire          rsp_xbar_demux_026_src0_valid;                                                                                          // rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_001:sink26_valid
	wire          rsp_xbar_demux_026_src0_startofpacket;                                                                                  // rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_001:sink26_startofpacket
	wire  [110:0] rsp_xbar_demux_026_src0_data;                                                                                           // rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_001:sink26_data
	wire   [37:0] rsp_xbar_demux_026_src0_channel;                                                                                        // rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_001:sink26_channel
	wire          rsp_xbar_demux_026_src0_ready;                                                                                          // rsp_xbar_mux_001:sink26_ready -> rsp_xbar_demux_026:src0_ready
	wire          rsp_xbar_demux_027_src0_endofpacket;                                                                                    // rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux_001:sink27_endofpacket
	wire          rsp_xbar_demux_027_src0_valid;                                                                                          // rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux_001:sink27_valid
	wire          rsp_xbar_demux_027_src0_startofpacket;                                                                                  // rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux_001:sink27_startofpacket
	wire  [110:0] rsp_xbar_demux_027_src0_data;                                                                                           // rsp_xbar_demux_027:src0_data -> rsp_xbar_mux_001:sink27_data
	wire   [37:0] rsp_xbar_demux_027_src0_channel;                                                                                        // rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux_001:sink27_channel
	wire          rsp_xbar_demux_027_src0_ready;                                                                                          // rsp_xbar_mux_001:sink27_ready -> rsp_xbar_demux_027:src0_ready
	wire          rsp_xbar_demux_029_src0_endofpacket;                                                                                    // rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux_001:sink29_endofpacket
	wire          rsp_xbar_demux_029_src0_valid;                                                                                          // rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux_001:sink29_valid
	wire          rsp_xbar_demux_029_src0_startofpacket;                                                                                  // rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux_001:sink29_startofpacket
	wire  [110:0] rsp_xbar_demux_029_src0_data;                                                                                           // rsp_xbar_demux_029:src0_data -> rsp_xbar_mux_001:sink29_data
	wire   [37:0] rsp_xbar_demux_029_src0_channel;                                                                                        // rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux_001:sink29_channel
	wire          rsp_xbar_demux_029_src0_ready;                                                                                          // rsp_xbar_mux_001:sink29_ready -> rsp_xbar_demux_029:src0_ready
	wire          rsp_xbar_demux_030_src0_endofpacket;                                                                                    // rsp_xbar_demux_030:src0_endofpacket -> rsp_xbar_mux_001:sink30_endofpacket
	wire          rsp_xbar_demux_030_src0_valid;                                                                                          // rsp_xbar_demux_030:src0_valid -> rsp_xbar_mux_001:sink30_valid
	wire          rsp_xbar_demux_030_src0_startofpacket;                                                                                  // rsp_xbar_demux_030:src0_startofpacket -> rsp_xbar_mux_001:sink30_startofpacket
	wire  [110:0] rsp_xbar_demux_030_src0_data;                                                                                           // rsp_xbar_demux_030:src0_data -> rsp_xbar_mux_001:sink30_data
	wire   [37:0] rsp_xbar_demux_030_src0_channel;                                                                                        // rsp_xbar_demux_030:src0_channel -> rsp_xbar_mux_001:sink30_channel
	wire          rsp_xbar_demux_030_src0_ready;                                                                                          // rsp_xbar_mux_001:sink30_ready -> rsp_xbar_demux_030:src0_ready
	wire          rsp_xbar_demux_032_src0_endofpacket;                                                                                    // rsp_xbar_demux_032:src0_endofpacket -> rsp_xbar_mux_001:sink32_endofpacket
	wire          rsp_xbar_demux_032_src0_valid;                                                                                          // rsp_xbar_demux_032:src0_valid -> rsp_xbar_mux_001:sink32_valid
	wire          rsp_xbar_demux_032_src0_startofpacket;                                                                                  // rsp_xbar_demux_032:src0_startofpacket -> rsp_xbar_mux_001:sink32_startofpacket
	wire  [110:0] rsp_xbar_demux_032_src0_data;                                                                                           // rsp_xbar_demux_032:src0_data -> rsp_xbar_mux_001:sink32_data
	wire   [37:0] rsp_xbar_demux_032_src0_channel;                                                                                        // rsp_xbar_demux_032:src0_channel -> rsp_xbar_mux_001:sink32_channel
	wire          rsp_xbar_demux_032_src0_ready;                                                                                          // rsp_xbar_mux_001:sink32_ready -> rsp_xbar_demux_032:src0_ready
	wire          rsp_xbar_demux_033_src0_endofpacket;                                                                                    // rsp_xbar_demux_033:src0_endofpacket -> rsp_xbar_mux_001:sink33_endofpacket
	wire          rsp_xbar_demux_033_src0_valid;                                                                                          // rsp_xbar_demux_033:src0_valid -> rsp_xbar_mux_001:sink33_valid
	wire          rsp_xbar_demux_033_src0_startofpacket;                                                                                  // rsp_xbar_demux_033:src0_startofpacket -> rsp_xbar_mux_001:sink33_startofpacket
	wire  [110:0] rsp_xbar_demux_033_src0_data;                                                                                           // rsp_xbar_demux_033:src0_data -> rsp_xbar_mux_001:sink33_data
	wire   [37:0] rsp_xbar_demux_033_src0_channel;                                                                                        // rsp_xbar_demux_033:src0_channel -> rsp_xbar_mux_001:sink33_channel
	wire          rsp_xbar_demux_033_src0_ready;                                                                                          // rsp_xbar_mux_001:sink33_ready -> rsp_xbar_demux_033:src0_ready
	wire          rsp_xbar_demux_034_src0_endofpacket;                                                                                    // rsp_xbar_demux_034:src0_endofpacket -> rsp_xbar_mux_001:sink34_endofpacket
	wire          rsp_xbar_demux_034_src0_valid;                                                                                          // rsp_xbar_demux_034:src0_valid -> rsp_xbar_mux_001:sink34_valid
	wire          rsp_xbar_demux_034_src0_startofpacket;                                                                                  // rsp_xbar_demux_034:src0_startofpacket -> rsp_xbar_mux_001:sink34_startofpacket
	wire  [110:0] rsp_xbar_demux_034_src0_data;                                                                                           // rsp_xbar_demux_034:src0_data -> rsp_xbar_mux_001:sink34_data
	wire   [37:0] rsp_xbar_demux_034_src0_channel;                                                                                        // rsp_xbar_demux_034:src0_channel -> rsp_xbar_mux_001:sink34_channel
	wire          rsp_xbar_demux_034_src0_ready;                                                                                          // rsp_xbar_mux_001:sink34_ready -> rsp_xbar_demux_034:src0_ready
	wire          rsp_xbar_demux_035_src0_endofpacket;                                                                                    // rsp_xbar_demux_035:src0_endofpacket -> rsp_xbar_mux_001:sink35_endofpacket
	wire          rsp_xbar_demux_035_src0_valid;                                                                                          // rsp_xbar_demux_035:src0_valid -> rsp_xbar_mux_001:sink35_valid
	wire          rsp_xbar_demux_035_src0_startofpacket;                                                                                  // rsp_xbar_demux_035:src0_startofpacket -> rsp_xbar_mux_001:sink35_startofpacket
	wire  [110:0] rsp_xbar_demux_035_src0_data;                                                                                           // rsp_xbar_demux_035:src0_data -> rsp_xbar_mux_001:sink35_data
	wire   [37:0] rsp_xbar_demux_035_src0_channel;                                                                                        // rsp_xbar_demux_035:src0_channel -> rsp_xbar_mux_001:sink35_channel
	wire          rsp_xbar_demux_035_src0_ready;                                                                                          // rsp_xbar_mux_001:sink35_ready -> rsp_xbar_demux_035:src0_ready
	wire          rsp_xbar_demux_036_src0_endofpacket;                                                                                    // rsp_xbar_demux_036:src0_endofpacket -> rsp_xbar_mux_001:sink36_endofpacket
	wire          rsp_xbar_demux_036_src0_valid;                                                                                          // rsp_xbar_demux_036:src0_valid -> rsp_xbar_mux_001:sink36_valid
	wire          rsp_xbar_demux_036_src0_startofpacket;                                                                                  // rsp_xbar_demux_036:src0_startofpacket -> rsp_xbar_mux_001:sink36_startofpacket
	wire  [110:0] rsp_xbar_demux_036_src0_data;                                                                                           // rsp_xbar_demux_036:src0_data -> rsp_xbar_mux_001:sink36_data
	wire   [37:0] rsp_xbar_demux_036_src0_channel;                                                                                        // rsp_xbar_demux_036:src0_channel -> rsp_xbar_mux_001:sink36_channel
	wire          rsp_xbar_demux_036_src0_ready;                                                                                          // rsp_xbar_mux_001:sink36_ready -> rsp_xbar_demux_036:src0_ready
	wire          rsp_xbar_demux_037_src0_endofpacket;                                                                                    // rsp_xbar_demux_037:src0_endofpacket -> rsp_xbar_mux_001:sink37_endofpacket
	wire          rsp_xbar_demux_037_src0_valid;                                                                                          // rsp_xbar_demux_037:src0_valid -> rsp_xbar_mux_001:sink37_valid
	wire          rsp_xbar_demux_037_src0_startofpacket;                                                                                  // rsp_xbar_demux_037:src0_startofpacket -> rsp_xbar_mux_001:sink37_startofpacket
	wire  [110:0] rsp_xbar_demux_037_src0_data;                                                                                           // rsp_xbar_demux_037:src0_data -> rsp_xbar_mux_001:sink37_data
	wire   [37:0] rsp_xbar_demux_037_src0_channel;                                                                                        // rsp_xbar_demux_037:src0_channel -> rsp_xbar_mux_001:sink37_channel
	wire          rsp_xbar_demux_037_src0_ready;                                                                                          // rsp_xbar_mux_001:sink37_ready -> rsp_xbar_demux_037:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                                            // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                                          // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [110:0] limiter_cmd_src_data;                                                                                                   // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [37:0] limiter_cmd_src_channel;                                                                                                // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                                  // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                           // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                                 // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                         // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [110:0] rsp_xbar_mux_src_data;                                                                                                  // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [37:0] rsp_xbar_mux_src_channel;                                                                                               // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                                 // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                                        // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                              // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                                      // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [110:0] addr_router_001_src_data;                                                                                               // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [37:0] addr_router_001_src_channel;                                                                                            // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                              // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                                       // rsp_xbar_mux_001:src_endofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                             // rsp_xbar_mux_001:src_valid -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                                     // rsp_xbar_mux_001:src_startofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [110:0] rsp_xbar_mux_001_src_data;                                                                                              // rsp_xbar_mux_001:src_data -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [37:0] rsp_xbar_mux_001_src_channel;                                                                                           // rsp_xbar_mux_001:src_channel -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                             // CPU_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                                        // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                              // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                                      // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [92:0] addr_router_002_src_data;                                                                                               // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [37:0] addr_router_002_src_channel;                                                                                            // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                              // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_016_src1_ready;                                                                                          // Video_In_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_016:src1_ready
	wire          addr_router_003_src_endofpacket;                                                                                        // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                                              // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                                      // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire   [92:0] addr_router_003_src_data;                                                                                               // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire   [37:0] addr_router_003_src_channel;                                                                                            // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                                              // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_demux_016_src2_ready;                                                                                          // Camera_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_016:src2_ready
	wire          addr_router_004_src_endofpacket;                                                                                        // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                                              // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                                      // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire   [92:0] addr_router_004_src_data;                                                                                               // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire   [37:0] addr_router_004_src_channel;                                                                                            // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                                              // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          rsp_xbar_demux_016_src3_ready;                                                                                          // LCD_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_016:src3_ready
	wire          addr_router_005_src_endofpacket;                                                                                        // addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          addr_router_005_src_valid;                                                                                              // addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	wire          addr_router_005_src_startofpacket;                                                                                      // addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire   [92:0] addr_router_005_src_data;                                                                                               // addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	wire   [37:0] addr_router_005_src_channel;                                                                                            // addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	wire          addr_router_005_src_ready;                                                                                              // cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	wire          rsp_xbar_demux_016_src4_ready;                                                                                          // VGA_DMA_Controller_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_016:src4_ready
	wire          addr_router_006_src_endofpacket;                                                                                        // addr_router_006:src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	wire          addr_router_006_src_valid;                                                                                              // addr_router_006:src_valid -> cmd_xbar_demux_006:sink_valid
	wire          addr_router_006_src_startofpacket;                                                                                      // addr_router_006:src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	wire   [92:0] addr_router_006_src_data;                                                                                               // addr_router_006:src_data -> cmd_xbar_demux_006:sink_data
	wire   [37:0] addr_router_006_src_channel;                                                                                            // addr_router_006:src_channel -> cmd_xbar_demux_006:sink_channel
	wire          addr_router_006_src_ready;                                                                                              // cmd_xbar_demux_006:sink_ready -> addr_router_006:src_ready
	wire          rsp_xbar_demux_016_src5_ready;                                                                                          // VideoConferencing_DMA_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_016:src5_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                           // cmd_xbar_mux:src_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                                 // cmd_xbar_mux:src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                         // cmd_xbar_mux:src_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_mux_src_data;                                                                                                  // cmd_xbar_mux:src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_mux_src_channel;                                                                                               // cmd_xbar_mux:src_channel -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                                 // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                              // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                                    // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                            // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [110:0] id_router_src_data;                                                                                                     // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [37:0] id_router_src_channel;                                                                                                  // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                                    // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                                       // cmd_xbar_mux_001:src_endofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                             // cmd_xbar_mux_001:src_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                                     // cmd_xbar_mux_001:src_startofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_mux_001_src_data;                                                                                              // cmd_xbar_mux_001:src_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_mux_001_src_channel;                                                                                           // cmd_xbar_mux_001:src_channel -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                             // SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                                          // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                                // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                        // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [110:0] id_router_001_src_data;                                                                                                 // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [37:0] id_router_001_src_channel;                                                                                              // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                                // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                                       // cmd_xbar_mux_002:src_endofpacket -> Flash_flash_data_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                             // cmd_xbar_mux_002:src_valid -> Flash_flash_data_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                                     // cmd_xbar_mux_002:src_startofpacket -> Flash_flash_data_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [110:0] cmd_xbar_mux_002_src_data;                                                                                              // cmd_xbar_mux_002:src_data -> Flash_flash_data_translator_avalon_universal_slave_0_agent:cp_data
	wire   [37:0] cmd_xbar_mux_002_src_channel;                                                                                           // cmd_xbar_mux_002:src_channel -> Flash_flash_data_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                             // Flash_flash_data_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                                          // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                                // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                                        // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [110:0] id_router_002_src_data;                                                                                                 // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [37:0] id_router_002_src_channel;                                                                                              // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                                // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                                          // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_003_src_endofpacket;                                                                                          // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                                // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                        // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [110:0] id_router_003_src_data;                                                                                                 // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [37:0] id_router_003_src_channel;                                                                                              // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                                // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                                          // Interval_Timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                                          // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                                // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                        // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [110:0] id_router_004_src_data;                                                                                                 // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [37:0] id_router_004_src_channel;                                                                                              // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                                // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                                          // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                                // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                                        // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [110:0] id_router_005_src_data;                                                                                                 // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [37:0] id_router_005_src_channel;                                                                                              // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                                // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                                          // Red_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                                          // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                                // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                        // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [110:0] id_router_006_src_data;                                                                                                 // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [37:0] id_router_006_src_channel;                                                                                              // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                                // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                                          // Green_LEDs_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                                          // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                                // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                        // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [110:0] id_router_007_src_data;                                                                                                 // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [37:0] id_router_007_src_channel;                                                                                              // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                                // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                                          // HEX3_HEX0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                                          // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                                // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                        // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [110:0] id_router_008_src_data;                                                                                                 // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [37:0] id_router_008_src_channel;                                                                                              // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                                // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                                          // HEX7_HEX4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_009_src_endofpacket;                                                                                          // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                                // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                        // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [110:0] id_router_009_src_data;                                                                                                 // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [37:0] id_router_009_src_channel;                                                                                              // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                                // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src10_ready;                                                                                         // Slider_Switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire          id_router_010_src_endofpacket;                                                                                          // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                                // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                                        // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [110:0] id_router_010_src_data;                                                                                                 // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [37:0] id_router_010_src_channel;                                                                                              // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                                // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_001_src11_ready;                                                                                         // Pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire          id_router_011_src_endofpacket;                                                                                          // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                                // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                                        // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [110:0] id_router_011_src_data;                                                                                                 // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [37:0] id_router_011_src_channel;                                                                                              // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                                // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                                         // Expansion_JP5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                                          // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                                // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                                        // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [110:0] id_router_012_src_data;                                                                                                 // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [37:0] id_router_012_src_channel;                                                                                              // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                                // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_001_src13_ready;                                                                                         // Serial_Port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire          id_router_013_src_endofpacket;                                                                                          // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                                // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                                        // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [110:0] id_router_013_src_data;                                                                                                 // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [37:0] id_router_013_src_channel;                                                                                              // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                                // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          width_adapter_src_ready;                                                                                                // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire          id_router_014_src_endofpacket;                                                                                          // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                                // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                                        // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire   [83:0] id_router_014_src_data;                                                                                                 // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [37:0] id_router_014_src_channel;                                                                                              // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                                // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_001_src15_ready;                                                                                         // PS2_Port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire          id_router_015_src_endofpacket;                                                                                          // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                                // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                                        // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [110:0] id_router_015_src_data;                                                                                                 // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [37:0] id_router_015_src_channel;                                                                                              // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                                // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_mux_016_src_endofpacket;                                                                                       // cmd_xbar_mux_016:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          cmd_xbar_mux_016_src_valid;                                                                                             // cmd_xbar_mux_016:src_valid -> burst_adapter_001:sink0_valid
	wire          cmd_xbar_mux_016_src_startofpacket;                                                                                     // cmd_xbar_mux_016:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [92:0] cmd_xbar_mux_016_src_data;                                                                                              // cmd_xbar_mux_016:src_data -> burst_adapter_001:sink0_data
	wire   [37:0] cmd_xbar_mux_016_src_channel;                                                                                           // cmd_xbar_mux_016:src_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_mux_016_src_ready;                                                                                             // burst_adapter_001:sink0_ready -> cmd_xbar_mux_016:src_ready
	wire          id_router_016_src_endofpacket;                                                                                          // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                                // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                                        // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire   [92:0] id_router_016_src_data;                                                                                                 // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [37:0] id_router_016_src_channel;                                                                                              // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                                // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_001_src17_ready;                                                                                         // VGA_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire          id_router_017_src_endofpacket;                                                                                          // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                                // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                                        // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [110:0] id_router_017_src_data;                                                                                                 // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [37:0] id_router_017_src_channel;                                                                                              // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                                // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          width_adapter_002_src_ready;                                                                                            // burst_adapter_002:sink0_ready -> width_adapter_002:out_ready
	wire          id_router_018_src_endofpacket;                                                                                          // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                                                // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                                        // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire   [83:0] id_router_018_src_data;                                                                                                 // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [37:0] id_router_018_src_channel;                                                                                              // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                                                // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_001_src19_ready;                                                                                         // OnBoard_AV_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src19_ready
	wire          id_router_019_src_endofpacket;                                                                                          // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                                                // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                                        // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [110:0] id_router_019_src_data;                                                                                                 // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [37:0] id_router_019_src_channel;                                                                                              // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                                                // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          cmd_xbar_demux_001_src20_ready;                                                                                         // PS2_Port_Dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src20_ready
	wire          id_router_020_src_endofpacket;                                                                                          // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                                                // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                                        // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [110:0] id_router_020_src_data;                                                                                                 // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [37:0] id_router_020_src_channel;                                                                                              // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                                                // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          cmd_xbar_demux_001_src21_ready;                                                                                         // Audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src21_ready
	wire          id_router_021_src_endofpacket;                                                                                          // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire          id_router_021_src_valid;                                                                                                // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire          id_router_021_src_startofpacket;                                                                                        // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [110:0] id_router_021_src_data;                                                                                                 // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire   [37:0] id_router_021_src_channel;                                                                                              // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire          id_router_021_src_ready;                                                                                                // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire          cmd_xbar_demux_001_src22_ready;                                                                                         // Flash_flash_erase_control_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src22_ready
	wire          id_router_022_src_endofpacket;                                                                                          // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire          id_router_022_src_valid;                                                                                                // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire          id_router_022_src_startofpacket;                                                                                        // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [110:0] id_router_022_src_data;                                                                                                 // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire   [37:0] id_router_022_src_channel;                                                                                              // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire          id_router_022_src_ready;                                                                                                // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire          cmd_xbar_demux_001_src23_ready;                                                                                         // SD_Card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src23_ready
	wire          id_router_023_src_endofpacket;                                                                                          // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire          id_router_023_src_valid;                                                                                                // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire          id_router_023_src_startofpacket;                                                                                        // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire  [110:0] id_router_023_src_data;                                                                                                 // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire   [37:0] id_router_023_src_channel;                                                                                              // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire          id_router_023_src_ready;                                                                                                // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire          cmd_xbar_demux_001_src24_ready;                                                                                         // IrDA_avalon_irda_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src24_ready
	wire          id_router_024_src_endofpacket;                                                                                          // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire          id_router_024_src_valid;                                                                                                // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire          id_router_024_src_startofpacket;                                                                                        // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire  [110:0] id_router_024_src_data;                                                                                                 // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire   [37:0] id_router_024_src_channel;                                                                                              // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire          id_router_024_src_ready;                                                                                                // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire          cmd_xbar_demux_001_src25_ready;                                                                                         // Video_In_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src25_ready
	wire          id_router_025_src_endofpacket;                                                                                          // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire          id_router_025_src_valid;                                                                                                // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire          id_router_025_src_startofpacket;                                                                                        // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire  [110:0] id_router_025_src_data;                                                                                                 // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire   [37:0] id_router_025_src_channel;                                                                                              // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire          id_router_025_src_ready;                                                                                                // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire          cmd_xbar_demux_001_src26_ready;                                                                                         // Camera_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src26_ready
	wire          id_router_026_src_endofpacket;                                                                                          // id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire          id_router_026_src_valid;                                                                                                // id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	wire          id_router_026_src_startofpacket;                                                                                        // id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire  [110:0] id_router_026_src_data;                                                                                                 // id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	wire   [37:0] id_router_026_src_channel;                                                                                              // id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	wire          id_router_026_src_ready;                                                                                                // rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	wire          cmd_xbar_demux_001_src27_ready;                                                                                         // Camera_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src27_ready
	wire          id_router_027_src_endofpacket;                                                                                          // id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire          id_router_027_src_valid;                                                                                                // id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	wire          id_router_027_src_startofpacket;                                                                                        // id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire  [110:0] id_router_027_src_data;                                                                                                 // id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	wire   [37:0] id_router_027_src_channel;                                                                                              // id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	wire          id_router_027_src_ready;                                                                                                // rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	wire          width_adapter_003_src_ready;                                                                                            // burst_adapter_003:sink0_ready -> width_adapter_003:out_ready
	wire          id_router_028_src_endofpacket;                                                                                          // id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire          id_router_028_src_valid;                                                                                                // id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	wire          id_router_028_src_startofpacket;                                                                                        // id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire   [83:0] id_router_028_src_data;                                                                                                 // id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	wire   [37:0] id_router_028_src_channel;                                                                                              // id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	wire          id_router_028_src_ready;                                                                                                // rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	wire          cmd_xbar_demux_001_src29_ready;                                                                                         // USB_avalon_usb_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src29_ready
	wire          id_router_029_src_endofpacket;                                                                                          // id_router_029:src_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	wire          id_router_029_src_valid;                                                                                                // id_router_029:src_valid -> rsp_xbar_demux_029:sink_valid
	wire          id_router_029_src_startofpacket;                                                                                        // id_router_029:src_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	wire  [110:0] id_router_029_src_data;                                                                                                 // id_router_029:src_data -> rsp_xbar_demux_029:sink_data
	wire   [37:0] id_router_029_src_channel;                                                                                              // id_router_029:src_channel -> rsp_xbar_demux_029:sink_channel
	wire          id_router_029_src_ready;                                                                                                // rsp_xbar_demux_029:sink_ready -> id_router_029:src_ready
	wire          cmd_xbar_demux_001_src30_ready;                                                                                         // LCD_Char_Buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src30_ready
	wire          id_router_030_src_endofpacket;                                                                                          // id_router_030:src_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	wire          id_router_030_src_valid;                                                                                                // id_router_030:src_valid -> rsp_xbar_demux_030:sink_valid
	wire          id_router_030_src_startofpacket;                                                                                        // id_router_030:src_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	wire  [110:0] id_router_030_src_data;                                                                                                 // id_router_030:src_data -> rsp_xbar_demux_030:sink_data
	wire   [37:0] id_router_030_src_channel;                                                                                              // id_router_030:src_channel -> rsp_xbar_demux_030:sink_channel
	wire          id_router_030_src_ready;                                                                                                // rsp_xbar_demux_030:sink_ready -> id_router_030:src_ready
	wire          width_adapter_004_src_ready;                                                                                            // burst_adapter_004:sink0_ready -> width_adapter_004:out_ready
	wire          id_router_031_src_endofpacket;                                                                                          // id_router_031:src_endofpacket -> rsp_xbar_demux_031:sink_endofpacket
	wire          id_router_031_src_valid;                                                                                                // id_router_031:src_valid -> rsp_xbar_demux_031:sink_valid
	wire          id_router_031_src_startofpacket;                                                                                        // id_router_031:src_startofpacket -> rsp_xbar_demux_031:sink_startofpacket
	wire   [83:0] id_router_031_src_data;                                                                                                 // id_router_031:src_data -> rsp_xbar_demux_031:sink_data
	wire   [37:0] id_router_031_src_channel;                                                                                              // id_router_031:src_channel -> rsp_xbar_demux_031:sink_channel
	wire          id_router_031_src_ready;                                                                                                // rsp_xbar_demux_031:sink_ready -> id_router_031:src_ready
	wire          cmd_xbar_demux_001_src32_ready;                                                                                         // enet_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src32_ready
	wire          id_router_032_src_endofpacket;                                                                                          // id_router_032:src_endofpacket -> rsp_xbar_demux_032:sink_endofpacket
	wire          id_router_032_src_valid;                                                                                                // id_router_032:src_valid -> rsp_xbar_demux_032:sink_valid
	wire          id_router_032_src_startofpacket;                                                                                        // id_router_032:src_startofpacket -> rsp_xbar_demux_032:sink_startofpacket
	wire  [110:0] id_router_032_src_data;                                                                                                 // id_router_032:src_data -> rsp_xbar_demux_032:sink_data
	wire   [37:0] id_router_032_src_channel;                                                                                              // id_router_032:src_channel -> rsp_xbar_demux_032:sink_channel
	wire          id_router_032_src_ready;                                                                                                // rsp_xbar_demux_032:sink_ready -> id_router_032:src_ready
	wire          cmd_xbar_demux_001_src33_ready;                                                                                         // packet_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src33_ready
	wire          id_router_033_src_endofpacket;                                                                                          // id_router_033:src_endofpacket -> rsp_xbar_demux_033:sink_endofpacket
	wire          id_router_033_src_valid;                                                                                                // id_router_033:src_valid -> rsp_xbar_demux_033:sink_valid
	wire          id_router_033_src_startofpacket;                                                                                        // id_router_033:src_startofpacket -> rsp_xbar_demux_033:sink_startofpacket
	wire  [110:0] id_router_033_src_data;                                                                                                 // id_router_033:src_data -> rsp_xbar_demux_033:sink_data
	wire   [37:0] id_router_033_src_channel;                                                                                              // id_router_033:src_channel -> rsp_xbar_demux_033:sink_channel
	wire          id_router_033_src_ready;                                                                                                // rsp_xbar_demux_033:sink_ready -> id_router_033:src_ready
	wire          cmd_xbar_demux_001_src34_ready;                                                                                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src34_ready
	wire          id_router_034_src_endofpacket;                                                                                          // id_router_034:src_endofpacket -> rsp_xbar_demux_034:sink_endofpacket
	wire          id_router_034_src_valid;                                                                                                // id_router_034:src_valid -> rsp_xbar_demux_034:sink_valid
	wire          id_router_034_src_startofpacket;                                                                                        // id_router_034:src_startofpacket -> rsp_xbar_demux_034:sink_startofpacket
	wire  [110:0] id_router_034_src_data;                                                                                                 // id_router_034:src_data -> rsp_xbar_demux_034:sink_data
	wire   [37:0] id_router_034_src_channel;                                                                                              // id_router_034:src_channel -> rsp_xbar_demux_034:sink_channel
	wire          id_router_034_src_ready;                                                                                                // rsp_xbar_demux_034:sink_ready -> id_router_034:src_ready
	wire          cmd_xbar_demux_001_src35_ready;                                                                                         // LCD_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src35_ready
	wire          id_router_035_src_endofpacket;                                                                                          // id_router_035:src_endofpacket -> rsp_xbar_demux_035:sink_endofpacket
	wire          id_router_035_src_valid;                                                                                                // id_router_035:src_valid -> rsp_xbar_demux_035:sink_valid
	wire          id_router_035_src_startofpacket;                                                                                        // id_router_035:src_startofpacket -> rsp_xbar_demux_035:sink_startofpacket
	wire  [110:0] id_router_035_src_data;                                                                                                 // id_router_035:src_data -> rsp_xbar_demux_035:sink_data
	wire   [37:0] id_router_035_src_channel;                                                                                              // id_router_035:src_channel -> rsp_xbar_demux_035:sink_channel
	wire          id_router_035_src_ready;                                                                                                // rsp_xbar_demux_035:sink_ready -> id_router_035:src_ready
	wire          cmd_xbar_demux_001_src36_ready;                                                                                         // VGA_DMA_Controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src36_ready
	wire          id_router_036_src_endofpacket;                                                                                          // id_router_036:src_endofpacket -> rsp_xbar_demux_036:sink_endofpacket
	wire          id_router_036_src_valid;                                                                                                // id_router_036:src_valid -> rsp_xbar_demux_036:sink_valid
	wire          id_router_036_src_startofpacket;                                                                                        // id_router_036:src_startofpacket -> rsp_xbar_demux_036:sink_startofpacket
	wire  [110:0] id_router_036_src_data;                                                                                                 // id_router_036:src_data -> rsp_xbar_demux_036:sink_data
	wire   [37:0] id_router_036_src_channel;                                                                                              // id_router_036:src_channel -> rsp_xbar_demux_036:sink_channel
	wire          id_router_036_src_ready;                                                                                                // rsp_xbar_demux_036:sink_ready -> id_router_036:src_ready
	wire          cmd_xbar_demux_001_src37_ready;                                                                                         // VideoConferencing_DMA_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src37_ready
	wire          id_router_037_src_endofpacket;                                                                                          // id_router_037:src_endofpacket -> rsp_xbar_demux_037:sink_endofpacket
	wire          id_router_037_src_valid;                                                                                                // id_router_037:src_valid -> rsp_xbar_demux_037:sink_valid
	wire          id_router_037_src_startofpacket;                                                                                        // id_router_037:src_startofpacket -> rsp_xbar_demux_037:sink_startofpacket
	wire  [110:0] id_router_037_src_data;                                                                                                 // id_router_037:src_data -> rsp_xbar_demux_037:sink_data
	wire   [37:0] id_router_037_src_channel;                                                                                              // id_router_037:src_channel -> rsp_xbar_demux_037:sink_channel
	wire          id_router_037_src_ready;                                                                                                // rsp_xbar_demux_037:sink_ready -> id_router_037:src_ready
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                                                   // cmd_xbar_demux_001:src14_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                                         // cmd_xbar_demux_001:src14_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                                                 // cmd_xbar_demux_001:src14_startofpacket -> width_adapter:in_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src14_data;                                                                                          // cmd_xbar_demux_001:src14_data -> width_adapter:in_data
	wire   [37:0] cmd_xbar_demux_001_src14_channel;                                                                                       // cmd_xbar_demux_001:src14_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_001_src14_ready;                                                                                         // width_adapter:in_ready -> cmd_xbar_demux_001:src14_ready
	wire          width_adapter_src_endofpacket;                                                                                          // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                                // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                                        // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [83:0] width_adapter_src_data;                                                                                                 // width_adapter:out_data -> burst_adapter:sink0_data
	wire   [37:0] width_adapter_src_channel;                                                                                              // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                                                   // cmd_xbar_demux_001:src16_endofpacket -> width_adapter_001:in_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                                         // cmd_xbar_demux_001:src16_valid -> width_adapter_001:in_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                                                 // cmd_xbar_demux_001:src16_startofpacket -> width_adapter_001:in_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src16_data;                                                                                          // cmd_xbar_demux_001:src16_data -> width_adapter_001:in_data
	wire   [37:0] cmd_xbar_demux_001_src16_channel;                                                                                       // cmd_xbar_demux_001:src16_channel -> width_adapter_001:in_channel
	wire          cmd_xbar_demux_001_src16_ready;                                                                                         // width_adapter_001:in_ready -> cmd_xbar_demux_001:src16_ready
	wire          width_adapter_001_src_endofpacket;                                                                                      // width_adapter_001:out_endofpacket -> cmd_xbar_mux_016:sink0_endofpacket
	wire          width_adapter_001_src_valid;                                                                                            // width_adapter_001:out_valid -> cmd_xbar_mux_016:sink0_valid
	wire          width_adapter_001_src_startofpacket;                                                                                    // width_adapter_001:out_startofpacket -> cmd_xbar_mux_016:sink0_startofpacket
	wire   [92:0] width_adapter_001_src_data;                                                                                             // width_adapter_001:out_data -> cmd_xbar_mux_016:sink0_data
	wire          width_adapter_001_src_ready;                                                                                            // cmd_xbar_mux_016:sink0_ready -> width_adapter_001:out_ready
	wire   [37:0] width_adapter_001_src_channel;                                                                                          // width_adapter_001:out_channel -> cmd_xbar_mux_016:sink0_channel
	wire          cmd_xbar_demux_001_src18_endofpacket;                                                                                   // cmd_xbar_demux_001:src18_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_001_src18_valid;                                                                                         // cmd_xbar_demux_001:src18_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_001_src18_startofpacket;                                                                                 // cmd_xbar_demux_001:src18_startofpacket -> width_adapter_002:in_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src18_data;                                                                                          // cmd_xbar_demux_001:src18_data -> width_adapter_002:in_data
	wire   [37:0] cmd_xbar_demux_001_src18_channel;                                                                                       // cmd_xbar_demux_001:src18_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_001_src18_ready;                                                                                         // width_adapter_002:in_ready -> cmd_xbar_demux_001:src18_ready
	wire          width_adapter_002_src_endofpacket;                                                                                      // width_adapter_002:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                                            // width_adapter_002:out_valid -> burst_adapter_002:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                                    // width_adapter_002:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire   [83:0] width_adapter_002_src_data;                                                                                             // width_adapter_002:out_data -> burst_adapter_002:sink0_data
	wire   [37:0] width_adapter_002_src_channel;                                                                                          // width_adapter_002:out_channel -> burst_adapter_002:sink0_channel
	wire          cmd_xbar_demux_001_src28_endofpacket;                                                                                   // cmd_xbar_demux_001:src28_endofpacket -> width_adapter_003:in_endofpacket
	wire          cmd_xbar_demux_001_src28_valid;                                                                                         // cmd_xbar_demux_001:src28_valid -> width_adapter_003:in_valid
	wire          cmd_xbar_demux_001_src28_startofpacket;                                                                                 // cmd_xbar_demux_001:src28_startofpacket -> width_adapter_003:in_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src28_data;                                                                                          // cmd_xbar_demux_001:src28_data -> width_adapter_003:in_data
	wire   [37:0] cmd_xbar_demux_001_src28_channel;                                                                                       // cmd_xbar_demux_001:src28_channel -> width_adapter_003:in_channel
	wire          cmd_xbar_demux_001_src28_ready;                                                                                         // width_adapter_003:in_ready -> cmd_xbar_demux_001:src28_ready
	wire          width_adapter_003_src_endofpacket;                                                                                      // width_adapter_003:out_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          width_adapter_003_src_valid;                                                                                            // width_adapter_003:out_valid -> burst_adapter_003:sink0_valid
	wire          width_adapter_003_src_startofpacket;                                                                                    // width_adapter_003:out_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire   [83:0] width_adapter_003_src_data;                                                                                             // width_adapter_003:out_data -> burst_adapter_003:sink0_data
	wire   [37:0] width_adapter_003_src_channel;                                                                                          // width_adapter_003:out_channel -> burst_adapter_003:sink0_channel
	wire          cmd_xbar_demux_001_src31_endofpacket;                                                                                   // cmd_xbar_demux_001:src31_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_001_src31_valid;                                                                                         // cmd_xbar_demux_001:src31_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_001_src31_startofpacket;                                                                                 // cmd_xbar_demux_001:src31_startofpacket -> width_adapter_004:in_startofpacket
	wire  [110:0] cmd_xbar_demux_001_src31_data;                                                                                          // cmd_xbar_demux_001:src31_data -> width_adapter_004:in_data
	wire   [37:0] cmd_xbar_demux_001_src31_channel;                                                                                       // cmd_xbar_demux_001:src31_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_001_src31_ready;                                                                                         // width_adapter_004:in_ready -> cmd_xbar_demux_001:src31_ready
	wire          width_adapter_004_src_endofpacket;                                                                                      // width_adapter_004:out_endofpacket -> burst_adapter_004:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                                                            // width_adapter_004:out_valid -> burst_adapter_004:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                                                    // width_adapter_004:out_startofpacket -> burst_adapter_004:sink0_startofpacket
	wire   [83:0] width_adapter_004_src_data;                                                                                             // width_adapter_004:out_data -> burst_adapter_004:sink0_data
	wire   [37:0] width_adapter_004_src_channel;                                                                                          // width_adapter_004:out_channel -> burst_adapter_004:sink0_channel
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                                    // rsp_xbar_demux_014:src0_endofpacket -> width_adapter_005:in_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                                          // rsp_xbar_demux_014:src0_valid -> width_adapter_005:in_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                                  // rsp_xbar_demux_014:src0_startofpacket -> width_adapter_005:in_startofpacket
	wire   [83:0] rsp_xbar_demux_014_src0_data;                                                                                           // rsp_xbar_demux_014:src0_data -> width_adapter_005:in_data
	wire   [37:0] rsp_xbar_demux_014_src0_channel;                                                                                        // rsp_xbar_demux_014:src0_channel -> width_adapter_005:in_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                                          // width_adapter_005:in_ready -> rsp_xbar_demux_014:src0_ready
	wire          width_adapter_005_src_endofpacket;                                                                                      // width_adapter_005:out_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          width_adapter_005_src_valid;                                                                                            // width_adapter_005:out_valid -> rsp_xbar_mux_001:sink14_valid
	wire          width_adapter_005_src_startofpacket;                                                                                    // width_adapter_005:out_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [110:0] width_adapter_005_src_data;                                                                                             // width_adapter_005:out_data -> rsp_xbar_mux_001:sink14_data
	wire          width_adapter_005_src_ready;                                                                                            // rsp_xbar_mux_001:sink14_ready -> width_adapter_005:out_ready
	wire   [37:0] width_adapter_005_src_channel;                                                                                          // width_adapter_005:out_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                                    // rsp_xbar_demux_016:src0_endofpacket -> width_adapter_006:in_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                                          // rsp_xbar_demux_016:src0_valid -> width_adapter_006:in_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                                  // rsp_xbar_demux_016:src0_startofpacket -> width_adapter_006:in_startofpacket
	wire   [92:0] rsp_xbar_demux_016_src0_data;                                                                                           // rsp_xbar_demux_016:src0_data -> width_adapter_006:in_data
	wire   [37:0] rsp_xbar_demux_016_src0_channel;                                                                                        // rsp_xbar_demux_016:src0_channel -> width_adapter_006:in_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                                          // width_adapter_006:in_ready -> rsp_xbar_demux_016:src0_ready
	wire          width_adapter_006_src_endofpacket;                                                                                      // width_adapter_006:out_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          width_adapter_006_src_valid;                                                                                            // width_adapter_006:out_valid -> rsp_xbar_mux_001:sink16_valid
	wire          width_adapter_006_src_startofpacket;                                                                                    // width_adapter_006:out_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [110:0] width_adapter_006_src_data;                                                                                             // width_adapter_006:out_data -> rsp_xbar_mux_001:sink16_data
	wire          width_adapter_006_src_ready;                                                                                            // rsp_xbar_mux_001:sink16_ready -> width_adapter_006:out_ready
	wire   [37:0] width_adapter_006_src_channel;                                                                                          // width_adapter_006:out_channel -> rsp_xbar_mux_001:sink16_channel
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                                    // rsp_xbar_demux_018:src0_endofpacket -> width_adapter_007:in_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                                          // rsp_xbar_demux_018:src0_valid -> width_adapter_007:in_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                                  // rsp_xbar_demux_018:src0_startofpacket -> width_adapter_007:in_startofpacket
	wire   [83:0] rsp_xbar_demux_018_src0_data;                                                                                           // rsp_xbar_demux_018:src0_data -> width_adapter_007:in_data
	wire   [37:0] rsp_xbar_demux_018_src0_channel;                                                                                        // rsp_xbar_demux_018:src0_channel -> width_adapter_007:in_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                                          // width_adapter_007:in_ready -> rsp_xbar_demux_018:src0_ready
	wire          width_adapter_007_src_endofpacket;                                                                                      // width_adapter_007:out_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire          width_adapter_007_src_valid;                                                                                            // width_adapter_007:out_valid -> rsp_xbar_mux_001:sink18_valid
	wire          width_adapter_007_src_startofpacket;                                                                                    // width_adapter_007:out_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [110:0] width_adapter_007_src_data;                                                                                             // width_adapter_007:out_data -> rsp_xbar_mux_001:sink18_data
	wire          width_adapter_007_src_ready;                                                                                            // rsp_xbar_mux_001:sink18_ready -> width_adapter_007:out_ready
	wire   [37:0] width_adapter_007_src_channel;                                                                                          // width_adapter_007:out_channel -> rsp_xbar_mux_001:sink18_channel
	wire          rsp_xbar_demux_028_src0_endofpacket;                                                                                    // rsp_xbar_demux_028:src0_endofpacket -> width_adapter_008:in_endofpacket
	wire          rsp_xbar_demux_028_src0_valid;                                                                                          // rsp_xbar_demux_028:src0_valid -> width_adapter_008:in_valid
	wire          rsp_xbar_demux_028_src0_startofpacket;                                                                                  // rsp_xbar_demux_028:src0_startofpacket -> width_adapter_008:in_startofpacket
	wire   [83:0] rsp_xbar_demux_028_src0_data;                                                                                           // rsp_xbar_demux_028:src0_data -> width_adapter_008:in_data
	wire   [37:0] rsp_xbar_demux_028_src0_channel;                                                                                        // rsp_xbar_demux_028:src0_channel -> width_adapter_008:in_channel
	wire          rsp_xbar_demux_028_src0_ready;                                                                                          // width_adapter_008:in_ready -> rsp_xbar_demux_028:src0_ready
	wire          width_adapter_008_src_endofpacket;                                                                                      // width_adapter_008:out_endofpacket -> rsp_xbar_mux_001:sink28_endofpacket
	wire          width_adapter_008_src_valid;                                                                                            // width_adapter_008:out_valid -> rsp_xbar_mux_001:sink28_valid
	wire          width_adapter_008_src_startofpacket;                                                                                    // width_adapter_008:out_startofpacket -> rsp_xbar_mux_001:sink28_startofpacket
	wire  [110:0] width_adapter_008_src_data;                                                                                             // width_adapter_008:out_data -> rsp_xbar_mux_001:sink28_data
	wire          width_adapter_008_src_ready;                                                                                            // rsp_xbar_mux_001:sink28_ready -> width_adapter_008:out_ready
	wire   [37:0] width_adapter_008_src_channel;                                                                                          // width_adapter_008:out_channel -> rsp_xbar_mux_001:sink28_channel
	wire          rsp_xbar_demux_031_src0_endofpacket;                                                                                    // rsp_xbar_demux_031:src0_endofpacket -> width_adapter_009:in_endofpacket
	wire          rsp_xbar_demux_031_src0_valid;                                                                                          // rsp_xbar_demux_031:src0_valid -> width_adapter_009:in_valid
	wire          rsp_xbar_demux_031_src0_startofpacket;                                                                                  // rsp_xbar_demux_031:src0_startofpacket -> width_adapter_009:in_startofpacket
	wire   [83:0] rsp_xbar_demux_031_src0_data;                                                                                           // rsp_xbar_demux_031:src0_data -> width_adapter_009:in_data
	wire   [37:0] rsp_xbar_demux_031_src0_channel;                                                                                        // rsp_xbar_demux_031:src0_channel -> width_adapter_009:in_channel
	wire          rsp_xbar_demux_031_src0_ready;                                                                                          // width_adapter_009:in_ready -> rsp_xbar_demux_031:src0_ready
	wire          width_adapter_009_src_endofpacket;                                                                                      // width_adapter_009:out_endofpacket -> rsp_xbar_mux_001:sink31_endofpacket
	wire          width_adapter_009_src_valid;                                                                                            // width_adapter_009:out_valid -> rsp_xbar_mux_001:sink31_valid
	wire          width_adapter_009_src_startofpacket;                                                                                    // width_adapter_009:out_startofpacket -> rsp_xbar_mux_001:sink31_startofpacket
	wire  [110:0] width_adapter_009_src_data;                                                                                             // width_adapter_009:out_data -> rsp_xbar_mux_001:sink31_data
	wire          width_adapter_009_src_ready;                                                                                            // rsp_xbar_mux_001:sink31_ready -> width_adapter_009:out_ready
	wire   [37:0] width_adapter_009_src_channel;                                                                                          // width_adapter_009:out_channel -> rsp_xbar_mux_001:sink31_channel
	wire   [37:0] limiter_cmd_valid_data;                                                                                                 // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                                               // JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                               // Interval_Timer:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                               // Serial_Port:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                               // Pushbuttons:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                                               // Expansion_JP5:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                                                               // PS2_Port:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                                                               // Audio:irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver7_irq;                                                                                               // PS2_Port_Dual:irq -> irq_mapper:receiver7_irq
	wire          irq_mapper_receiver8_irq;                                                                                               // IrDA:irq -> irq_mapper:receiver8_irq
	wire          irq_mapper_receiver9_irq;                                                                                               // Accelerometer:irq -> irq_mapper:receiver9_irq
	wire          irq_mapper_receiver10_irq;                                                                                              // USB:irq -> irq_mapper:receiver10_irq
	wire          irq_mapper_receiver11_irq;                                                                                              // Slider_Switches:irq -> irq_mapper:receiver11_irq
	wire   [31:0] cpu_d_irq_irq;                                                                                                          // irq_mapper:sender_irq -> CPU:d_irq
	wire          enet_receive_endofpacket;                                                                                               // enet:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire          enet_receive_valid;                                                                                                     // enet:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire          enet_receive_startofpacket;                                                                                             // enet:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire    [5:0] enet_receive_error;                                                                                                     // enet:rx_err -> avalon_st_adapter:in_0_error
	wire    [1:0] enet_receive_empty;                                                                                                     // enet:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire   [31:0] enet_receive_data;                                                                                                      // enet:ff_rx_data -> avalon_st_adapter:in_0_data
	wire          enet_receive_ready;                                                                                                     // avalon_st_adapter:in_0_ready -> enet:ff_rx_rdy
	wire          avalon_st_adapter_out_0_endofpacket;                                                                                    // avalon_st_adapter:out_0_endofpacket -> VideoConferencing_DMA_0:eth_rx_eop
	wire          avalon_st_adapter_out_0_valid;                                                                                          // avalon_st_adapter:out_0_valid -> VideoConferencing_DMA_0:eth_rx_dval
	wire          avalon_st_adapter_out_0_startofpacket;                                                                                  // avalon_st_adapter:out_0_startofpacket -> VideoConferencing_DMA_0:eth_rx_sop
	wire    [5:0] avalon_st_adapter_out_0_error;                                                                                          // avalon_st_adapter:out_0_error -> VideoConferencing_DMA_0:eth_rx_error
	wire   [31:0] avalon_st_adapter_out_0_data;                                                                                           // avalon_st_adapter:out_0_data -> VideoConferencing_DMA_0:eth_rx_data
	wire    [1:0] avalon_st_adapter_out_0_channel;                                                                                        // avalon_st_adapter:out_0_channel -> VideoConferencing_DMA_0:eth_rx_mod
	wire          avalon_st_adapter_out_0_ready;                                                                                          // VideoConferencing_DMA_0:eth_rx_rdy -> avalon_st_adapter:out_0_ready
	wire          videoconferencing_dma_0_avalon_streaming_source_endofpacket;                                                            // VideoConferencing_DMA_0:eth_tx_eop -> avalon_st_adapter_001:in_0_endofpacket
	wire          videoconferencing_dma_0_avalon_streaming_source_valid;                                                                  // VideoConferencing_DMA_0:eth_tx_wren -> avalon_st_adapter_001:in_0_valid
	wire          videoconferencing_dma_0_avalon_streaming_source_startofpacket;                                                          // VideoConferencing_DMA_0:eth_tx_sop -> avalon_st_adapter_001:in_0_startofpacket
	wire    [5:0] videoconferencing_dma_0_avalon_streaming_source_error;                                                                  // VideoConferencing_DMA_0:eth_tx_error -> avalon_st_adapter_001:in_0_error
	wire   [31:0] videoconferencing_dma_0_avalon_streaming_source_data;                                                                   // VideoConferencing_DMA_0:eth_tx_data -> avalon_st_adapter_001:in_0_data
	wire    [1:0] videoconferencing_dma_0_avalon_streaming_source_channel;                                                                // VideoConferencing_DMA_0:eth_tx_mod -> avalon_st_adapter_001:in_0_channel
	wire          videoconferencing_dma_0_avalon_streaming_source_ready;                                                                  // avalon_st_adapter_001:in_0_ready -> VideoConferencing_DMA_0:eth_tx_rdy
	wire          avalon_st_adapter_001_out_0_endofpacket;                                                                                // avalon_st_adapter_001:out_0_endofpacket -> enet:ff_tx_eop
	wire          avalon_st_adapter_001_out_0_valid;                                                                                      // avalon_st_adapter_001:out_0_valid -> enet:ff_tx_wren
	wire          avalon_st_adapter_001_out_0_startofpacket;                                                                              // avalon_st_adapter_001:out_0_startofpacket -> enet:ff_tx_sop
	wire    [0:0] avalon_st_adapter_001_out_0_error;                                                                                      // avalon_st_adapter_001:out_0_error -> enet:ff_tx_err
	wire    [1:0] avalon_st_adapter_001_out_0_empty;                                                                                      // avalon_st_adapter_001:out_0_empty -> enet:ff_tx_mod
	wire   [31:0] avalon_st_adapter_001_out_0_data;                                                                                       // avalon_st_adapter_001:out_0_data -> enet:ff_tx_data
	wire          avalon_st_adapter_001_out_0_ready;                                                                                      // enet:ff_tx_rdy -> avalon_st_adapter_001:out_0_ready

	nios_system_JTAG_UART jtag_uart (
		.clk            (sys_clk),                                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	nios_system_Interval_Timer interval_timer (
		.clk        (sys_clk),                                                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                             // reset.reset_n
		.address    (interval_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (interval_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (interval_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (interval_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~interval_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                                     //   irq.irq
	);

	nios_system_SDRAM sdram (
		.clk            (sys_clk),                                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                       // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_SDRAM),                                //  wire.export
		.zs_ba          (zs_ba_from_the_SDRAM),                                  //      .export
		.zs_cas_n       (zs_cas_n_from_the_SDRAM),                               //      .export
		.zs_cke         (zs_cke_from_the_SDRAM),                                 //      .export
		.zs_cs_n        (zs_cs_n_from_the_SDRAM),                                //      .export
		.zs_dq          (zs_dq_to_and_from_the_SDRAM),                           //      .export
		.zs_dqm         (zs_dqm_from_the_SDRAM),                                 //      .export
		.zs_ras_n       (zs_ras_n_from_the_SDRAM),                               //      .export
		.zs_we_n        (zs_we_n_from_the_SDRAM)                                 //      .export
	);

	nios_system_Red_LEDs red_leds (
		.clk        (sys_clk),                                                                       //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                //          clock_reset_reset.reset
		.address    (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.LEDR       (LEDR_from_the_Red_LEDs)                                                         //         external_interface.export
	);

	nios_system_Green_LEDs green_leds (
		.clk        (sys_clk),                                                                         //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                  //          clock_reset_reset.reset
		.address    (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.LEDG       (LEDG_from_the_Green_LEDs)                                                         //         external_interface.export
	);

	nios_system_HEX3_HEX0 hex3_hex0 (
		.clk        (sys_clk),                                                                        //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                 //          clock_reset_reset.reset
		.address    (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.HEX0       (HEX0_from_the_HEX3_HEX0),                                                        //         external_interface.export
		.HEX1       (HEX1_from_the_HEX3_HEX0),                                                        //                           .export
		.HEX2       (HEX2_from_the_HEX3_HEX0),                                                        //                           .export
		.HEX3       (HEX3_from_the_HEX3_HEX0)                                                         //                           .export
	);

	nios_system_HEX7_HEX4 hex7_hex4 (
		.clk        (sys_clk),                                                                        //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                 //          clock_reset_reset.reset
		.address    (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.HEX4       (HEX4_from_the_HEX7_HEX4),                                                        //         external_interface.export
		.HEX5       (HEX5_from_the_HEX7_HEX4),                                                        //                           .export
		.HEX6       (HEX6_from_the_HEX7_HEX4),                                                        //                           .export
		.HEX7       (HEX7_from_the_HEX7_HEX4)                                                         //                           .export
	);

	nios_system_Slider_Switches slider_switches (
		.clk        (sys_clk),                                                                              //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                       //          clock_reset_reset.reset
		.address    (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.in_port    (Slider_Switches_external_interface_export),                                            //         external_interface.export
		.irq        (irq_mapper_receiver11_irq)                                                             //                  interrupt.irq
	);

	nios_system_Pushbuttons pushbuttons (
		.clk        (sys_clk),                                                                          //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                   //          clock_reset_reset.reset
		.address    (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.KEY        (KEY_to_the_Pushbuttons),                                                           //         external_interface.export
		.irq        (irq_mapper_receiver3_irq)                                                          //                  interrupt.irq
	);

	nios_system_Expansion_JP5 expansion_jp5 (
		.clk        (sys_clk),                                                                            //                clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                                     //          clock_reset_reset.reset
		.address    (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),    // avalon_parallel_port_slave.address
		.byteenable (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.chipselect (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.read       (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.write      (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.writedata  (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.readdata   (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.GPIO       (GPIO_to_and_from_the_Expansion_JP5),                                                 //         external_interface.export
		.irq        (irq_mapper_receiver4_irq)                                                            //                  interrupt.irq
	);

	nios_system_Serial_Port serial_port (
		.clk        (sys_clk),                                                                  //        clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                           //  clock_reset_reset.reset
		.address    (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_address),    // avalon_rs232_slave.address
		.chipselect (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.byteenable (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable), //                   .byteenable
		.read       (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write      (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata  (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata   (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver2_irq),                                                 //          interrupt.irq
		.UART_RXD   (UART_RXD_to_the_Serial_Port),                                              // external_interface.export
		.UART_TXD   (UART_TXD_from_the_Serial_Port)                                             //                   .export
	);

	nios_system_OnBoard_AV onboard_av (
		.clk         (sys_clk),                                                                      //            clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                               //      clock_reset_reset.reset
		.address     (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_address),     // avalon_av_config_slave.address
		.byteenable  (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),  //                       .byteenable
		.read        (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_read),        //                       .read
		.write       (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_write),       //                       .write
		.writedata   (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),   //                       .writedata
		.readdata    (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),    //                       .readdata
		.waitrequest (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest), //                       .waitrequest
		.I2C_SDAT    (I2C_SDAT_to_and_from_the_AV_Config),                                           //     external_interface.export
		.I2C_SCLK    (I2C_SCLK_from_the_AV_Config)                                                   //                       .export
	);

	nios_system_Audio audio (
		.clk         (sys_clk),                                                            //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                     //  clock_reset_reset.reset
		.address     (audio_avalon_audio_slave_translator_avalon_anti_slave_0_address),    // avalon_audio_slave.address
		.chipselect  (audio_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.read        (audio_avalon_audio_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write       (audio_avalon_audio_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata   (audio_avalon_audio_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata    (audio_avalon_audio_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver6_irq),                                           //          interrupt.irq
		.AUD_ADCDAT  (AUD_ADCDAT_to_the_Audio),                                            // external_interface.export
		.AUD_ADCLRCK (AUD_ADCLRCK_to_the_Audio),                                           //                   .export
		.AUD_BCLK    (AUD_BCLK_to_the_Audio),                                              //                   .export
		.AUD_DACDAT  (AUD_DACDAT_from_the_Audio),                                          //                   .export
		.AUD_DACLRCK (AUD_DACLRCK_to_the_Audio)                                            //                   .export
	);

	nios_system_Char_LCD_16x2 char_lcd_16x2 (
		.clk         (sys_clk),                                                                   //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                            //  clock_reset_reset.reset
		.address     (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_address),     //   avalon_lcd_slave.address
		.chipselect  (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.read        (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.LCD_DATA    (LCD_DATA_to_and_from_the_Char_LCD_16x2),                                    // external_interface.export
		.LCD_ON      (LCD_ON_from_the_Char_LCD_16x2),                                             //                   .export
		.LCD_BLON    (LCD_BLON_from_the_Char_LCD_16x2),                                           //                   .export
		.LCD_EN      (LCD_EN_from_the_Char_LCD_16x2),                                             //                   .export
		.LCD_RS      (LCD_RS_from_the_Char_LCD_16x2),                                             //                   .export
		.LCD_RW      (LCD_RW_from_the_Char_LCD_16x2)                                              //                   .export
	);

	nios_system_PS2_Port ps2_port (
		.clk         (sys_clk),                                                              //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                       //  clock_reset_reset.reset
		.address     (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_address),     //   avalon_ps2_slave.address
		.chipselect  (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.byteenable  (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable),  //                   .byteenable
		.read        (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver5_irq),                                             //          interrupt.irq
		.PS2_CLK     (PS2_CLK_to_and_from_the_PS2_Port),                                     // external_interface.export
		.PS2_DAT     (PS2_DAT_to_and_from_the_PS2_Port)                                      //                   .export
	);

	nios_system_SRAM sram (
		.clk           (sys_clk),                                                             //        clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                      //  clock_reset_reset.reset
		.SRAM_DQ       (SRAM_DQ_to_and_from_the_SRAM),                                        // external_interface.export
		.SRAM_ADDR     (SRAM_ADDR_from_the_SRAM),                                             //                   .export
		.SRAM_LB_N     (SRAM_LB_N_from_the_SRAM),                                             //                   .export
		.SRAM_UB_N     (SRAM_UB_N_from_the_SRAM),                                             //                   .export
		.SRAM_CE_N     (SRAM_CE_N_from_the_SRAM),                                             //                   .export
		.SRAM_OE_N     (SRAM_OE_N_from_the_SRAM),                                             //                   .export
		.SRAM_WE_N     (SRAM_WE_N_from_the_SRAM),                                             //                   .export
		.address       (sram_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (sram_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (sram_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	nios_system_VGA_Char_Buffer vga_char_buffer (
		.clk                  (sys_clk),                                                                             //               clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                      //         clock_reset_reset.reset
		.ctrl_address         (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable), //                          .byteenable
		.ctrl_chipselect      (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect), //                          .chipselect
		.ctrl_read            (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read),       //                          .read
		.ctrl_write           (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write),      //                          .write
		.ctrl_writedata       (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),  //                          .writedata
		.ctrl_readdata        (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),   //                          .readdata
		.buf_byteenable       (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),  //                          .chipselect
		.buf_read             (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),        //                          .read
		.buf_write            (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),       //                          .write
		.buf_writedata        (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.buf_readdata         (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.buf_waitrequest      (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.buf_address          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),     //                          .address
		.stream_ready         (vga_char_buffer_avalon_char_source_ready),                                            //        avalon_char_source.ready
		.stream_startofpacket (vga_char_buffer_avalon_char_source_startofpacket),                                    //                          .startofpacket
		.stream_endofpacket   (vga_char_buffer_avalon_char_source_endofpacket),                                      //                          .endofpacket
		.stream_valid         (vga_char_buffer_avalon_char_source_valid),                                            //                          .valid
		.stream_data          (vga_char_buffer_avalon_char_source_data)                                              //                          .data
	);

	nios_system_VGA_Controller vga_controller (
		.clk           (vga_clk_out_clk_clk),                                       //        clock_reset.clk
		.reset         (rst_controller_001_reset_out_reset),                        //  clock_reset_reset.reset
		.data          (vga_dual_clock_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (vga_dual_clock_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (vga_dual_clock_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_external_interface_CLK),                     // external_interface.export
		.VGA_HS        (vga_controller_external_interface_HS),                      //                   .export
		.VGA_VS        (vga_controller_external_interface_VS),                      //                   .export
		.VGA_BLANK     (vga_controller_external_interface_BLANK),                   //                   .export
		.VGA_SYNC      (vga_controller_external_interface_SYNC),                    //                   .export
		.VGA_R         (vga_controller_external_interface_R),                       //                   .export
		.VGA_G         (vga_controller_external_interface_G),                       //                   .export
		.VGA_B         (vga_controller_external_interface_B)                        //                   .export
	);

	nios_system_VGA_Pixel_RGB_Resampler vga_pixel_rgb_resampler (
		.clk                      (sys_clk),                                                 //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                          // clock_reset_reset.reset
		.stream_in_startofpacket  (vga_dma_controller_avalon_pixel_source_startofpacket),    //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (vga_dma_controller_avalon_pixel_source_endofpacket),      //                  .endofpacket
		.stream_in_valid          (vga_dma_controller_avalon_pixel_source_valid),            //                  .valid
		.stream_in_ready          (vga_dma_controller_avalon_pixel_source_ready),            //                  .ready
		.stream_in_data           (vga_dma_controller_avalon_pixel_source_data),             //                  .data
		.stream_out_ready         (vga_pixel_rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (vga_pixel_rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (vga_pixel_rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	nios_system_VGA_Pixel_Scaler vga_pixel_scaler (
		.clk                      (sys_clk),                                                 //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                          //    clock_reset_reset.reset
		.stream_in_startofpacket  (vga_pixel_rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (vga_pixel_rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (vga_pixel_rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (vga_pixel_rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (vga_pixel_rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (vga_pixel_scaler_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (vga_pixel_scaler_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (vga_pixel_scaler_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (vga_pixel_scaler_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (vga_pixel_scaler_avalon_scaler_source_data)               //                     .data
	);

	nios_system_VGA_Dual_Clock_FIFO vga_dual_clock_fifo (
		.clk_stream_in            (sys_clk),                                                   //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                            //   clock_stream_in_reset.reset
		.clk_stream_out           (vga_clk_out_clk_clk),                                       //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_001_reset_out_reset),                        //  clock_stream_out_reset.reset
		.stream_in_ready          (vga_alpha_blender_avalon_blended_source_ready),             //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (vga_alpha_blender_avalon_blended_source_startofpacket),     //                        .startofpacket
		.stream_in_endofpacket    (vga_alpha_blender_avalon_blended_source_endofpacket),       //                        .endofpacket
		.stream_in_valid          (vga_alpha_blender_avalon_blended_source_valid),             //                        .valid
		.stream_in_data           (vga_alpha_blender_avalon_blended_source_data),              //                        .data
		.stream_out_ready         (vga_dual_clock_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (vga_dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (vga_dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (vga_dual_clock_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (vga_dual_clock_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	fpoint_wrapper #(
		.useDivider (1)
	) cpu_fpoint (
		.clk    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk),    // s1.clk
		.clk_en (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //   .clk_en
		.dataa  (cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //   .dataa
		.datab  (cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //   .datab
		.n      (cpu_custom_instruction_master_multi_slave_translator0_ci_master_n),      //   .n
		.reset  (cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //   .reset
		.start  (cpu_custom_instruction_master_multi_slave_translator0_ci_master_start),  //   .start
		.done   (cpu_custom_instruction_master_multi_slave_translator0_ci_master_done),   //   .done
		.result (cpu_custom_instruction_master_multi_slave_translator0_ci_master_result)  //   .result
	);

	nios_system_VGA_Alpha_Blender vga_alpha_blender (
		.clk                      (sys_clk),                                               //            clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                        //      clock_reset_reset.reset
		.foreground_data          (vga_char_buffer_avalon_char_source_data),               // avalon_foreground_sink.data
		.foreground_startofpacket (vga_char_buffer_avalon_char_source_startofpacket),      //                       .startofpacket
		.foreground_endofpacket   (vga_char_buffer_avalon_char_source_endofpacket),        //                       .endofpacket
		.foreground_valid         (vga_char_buffer_avalon_char_source_valid),              //                       .valid
		.foreground_ready         (vga_char_buffer_avalon_char_source_ready),              //                       .ready
		.background_data          (vga_pixel_scaler_avalon_scaler_source_data),            // avalon_background_sink.data
		.background_startofpacket (vga_pixel_scaler_avalon_scaler_source_startofpacket),   //                       .startofpacket
		.background_endofpacket   (vga_pixel_scaler_avalon_scaler_source_endofpacket),     //                       .endofpacket
		.background_valid         (vga_pixel_scaler_avalon_scaler_source_valid),           //                       .valid
		.background_ready         (vga_pixel_scaler_avalon_scaler_source_ready),           //                       .ready
		.output_ready             (vga_alpha_blender_avalon_blended_source_ready),         //  avalon_blended_source.ready
		.output_data              (vga_alpha_blender_avalon_blended_source_data),          //                       .data
		.output_startofpacket     (vga_alpha_blender_avalon_blended_source_startofpacket), //                       .startofpacket
		.output_endofpacket       (vga_alpha_blender_avalon_blended_source_endofpacket),   //                       .endofpacket
		.output_valid             (vga_alpha_blender_avalon_blended_source_valid)          //                       .valid
	);

	nios_system_PS2_Port ps2_port_dual (
		.clk         (sys_clk),                                                                   //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                            //  clock_reset_reset.reset
		.address     (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_address),     //   avalon_ps2_slave.address
		.chipselect  (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.byteenable  (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable),  //                   .byteenable
		.read        (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver7_irq),                                                  //          interrupt.irq
		.PS2_CLK     (PS2_CLK_to_and_from_the_PS2_Port_Dual),                                     // external_interface.export
		.PS2_DAT     (PS2_DAT_to_and_from_the_PS2_Port_Dual)                                      //                   .export
	);

	nios_system_CPU cpu (
		.clk                                   (sys_clk),                                                          //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                  //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                          //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (cpu_data_master_read),                                             //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                            //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                      //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.A_ci_multi_done                       (cpu_custom_instruction_master_done),                               // custom_instruction_master.done
		.A_ci_multi_result                     (cpu_custom_instruction_master_multi_result),                       //                          .multi_result
		.A_ci_multi_a                          (cpu_custom_instruction_master_multi_a),                            //                          .multi_a
		.A_ci_multi_b                          (cpu_custom_instruction_master_multi_b),                            //                          .multi_b
		.A_ci_multi_c                          (cpu_custom_instruction_master_multi_c),                            //                          .multi_c
		.A_ci_multi_clk_en                     (cpu_custom_instruction_master_clk_en),                             //                          .clk_en
		.A_ci_multi_clock                      (cpu_custom_instruction_master_clk),                                //                          .clk
		.A_ci_multi_reset                      (cpu_custom_instruction_master_reset),                              //                          .reset
		.A_ci_multi_dataa                      (cpu_custom_instruction_master_multi_dataa),                        //                          .multi_dataa
		.A_ci_multi_datab                      (cpu_custom_instruction_master_multi_datab),                        //                          .multi_datab
		.A_ci_multi_n                          (cpu_custom_instruction_master_multi_n),                            //                          .multi_n
		.A_ci_multi_readra                     (cpu_custom_instruction_master_multi_readra),                       //                          .multi_readra
		.A_ci_multi_readrb                     (cpu_custom_instruction_master_multi_readrb),                       //                          .multi_readrb
		.A_ci_multi_start                      (cpu_custom_instruction_master_start),                              //                          .start
		.A_ci_multi_writerc                    (cpu_custom_instruction_master_multi_writerc)                       //                          .multi_writerc
	);

	nios_system_sysid sysid (
		.clock    (sys_clk),                                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                             //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	nios_system_External_Clocks external_clocks (
		.CLOCK_50    (clk),                                //       clk_in_primary.clk
		.reset       (rst_controller_002_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (sys_clk),                            //              sys_clk.clk
		.sys_reset_n (),                                   //        sys_clk_reset.reset_n
		.SDRAM_CLK   (sdram_clk),                          //            sdram_clk.clk
		.VGA_CLK     (vga_clk_out_clk_clk),                //              vga_clk.clk
		.VGA_CLK_33  (external_clocks_vga_clk_33_clk),     //           vga_clk_33.clk
		.CLOCK_27    (clk_27),                             //     clk_in_secondary.clk
		.AUD_CLK     (audio_clk)                           //            audio_clk.clk
	);

	Altera_UP_Flash_Memory_IP_Core_Avalon_Interface flash (
		.i_avalon_chip_select       (flash_flash_data_translator_avalon_anti_slave_0_chipselect),           //          flash_data.chipselect
		.i_avalon_write             (flash_flash_data_translator_avalon_anti_slave_0_write),                //                    .write
		.i_avalon_read              (flash_flash_data_translator_avalon_anti_slave_0_read),                 //                    .read
		.i_avalon_address           (flash_flash_data_translator_avalon_anti_slave_0_address),              //                    .address
		.i_avalon_byteenable        (flash_flash_data_translator_avalon_anti_slave_0_byteenable),           //                    .byteenable
		.i_avalon_writedata         (flash_flash_data_translator_avalon_anti_slave_0_writedata),            //                    .writedata
		.o_avalon_readdata          (flash_flash_data_translator_avalon_anti_slave_0_readdata),             //                    .readdata
		.o_avalon_waitrequest       (flash_flash_data_translator_avalon_anti_slave_0_waitrequest),          //                    .waitrequest
		.i_clock                    (sys_clk),                                                              //          clock_sink.clk
		.i_reset_n                  (~rst_controller_003_reset_out_reset),                                  //    clock_sink_reset.reset_n
		.FL_ADDR                    (flash_ADDR),                                                           //         conduit_end.export
		.FL_CE_N                    (flash_CE_N),                                                           //                    .export
		.FL_OE_N                    (flash_OE_N),                                                           //                    .export
		.FL_WE_N                    (flash_WE_N),                                                           //                    .export
		.FL_RST_N                   (flash_RST_N),                                                          //                    .export
		.FL_DQ                      (flash_DQ),                                                             //                    .export
		.i_avalon_erase_write       (flash_flash_erase_control_translator_avalon_anti_slave_0_write),       // flash_erase_control.write
		.i_avalon_erase_read        (flash_flash_erase_control_translator_avalon_anti_slave_0_read),        //                    .read
		.i_avalon_erase_byteenable  (flash_flash_erase_control_translator_avalon_anti_slave_0_byteenable),  //                    .byteenable
		.i_avalon_erase_writedata   (flash_flash_erase_control_translator_avalon_anti_slave_0_writedata),   //                    .writedata
		.i_avalon_erase_chip_select (flash_flash_erase_control_translator_avalon_anti_slave_0_chipselect),  //                    .chipselect
		.o_avalon_erase_readdata    (flash_flash_erase_control_translator_avalon_anti_slave_0_readdata),    //                    .readdata
		.o_avalon_erase_waitrequest (flash_flash_erase_control_translator_avalon_anti_slave_0_waitrequest)  //                    .waitrequest
	);

	Altera_UP_SD_Card_Avalon_Interface sd_card (
		.i_avalon_chip_select (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),     //                    .address
		.i_avalon_read        (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),        //                    .read
		.i_avalon_write       (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),       //                    .write
		.i_avalon_byteenable  (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),  //                    .byteenable
		.i_avalon_writedata   (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),   //                    .writedata
		.o_avalon_readdata    (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),    //                    .readdata
		.o_avalon_waitrequest (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest), //                    .waitrequest
		.i_clock              (sys_clk),                                                                //          clock_sink.clk
		.i_reset_n            (~rst_controller_003_reset_out_reset),                                    //    clock_sink_reset.reset_n
		.b_SD_cmd             (sdcard_b_SD_cmd),                                                        //         conduit_end.export
		.b_SD_dat             (sdcard_b_SD_dat),                                                        //                    .export
		.b_SD_dat3            (sdcard_b_SD_dat3),                                                       //                    .export
		.o_SD_clock           (sdcard_o_SD_clock)                                                       //                    .export
	);

	nios_system_IrDA irda (
		.clk        (sys_clk),                                                          //        clock_reset.clk
		.reset      (rst_controller_003_reset_out_reset),                               //  clock_reset_reset.reset
		.address    (irda_avalon_irda_slave_translator_avalon_anti_slave_0_address),    //  avalon_irda_slave.address
		.chipselect (irda_avalon_irda_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.byteenable (irda_avalon_irda_slave_translator_avalon_anti_slave_0_byteenable), //                   .byteenable
		.read       (irda_avalon_irda_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write      (irda_avalon_irda_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata  (irda_avalon_irda_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata   (irda_avalon_irda_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver8_irq),                                         //          interrupt.irq
		.IRDA_TXD   (irda_TXD),                                                         // external_interface.export
		.IRDA_RXD   (irda_RXD)                                                          //                   .export
	);

	nios_system_Video_In video_in (
		.clk                      (sys_clk),                                      //           clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),               //     clock_reset_reset.reset
		.stream_out_ready         (video_in_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (video_in_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (video_in_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (video_in_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (video_in_avalon_decoder_source_data),          //                      .data
		.TD_CLK27                 (video_in_TD_CLK27),                            //    external_interface.export
		.TD_DATA                  (video_in_TD_DATA),                             //                      .export
		.TD_HS                    (video_in_TD_HS),                               //                      .export
		.TD_VS                    (video_in_TD_VS),                               //                      .export
		.clk27_reset              (video_in_clk27_reset),                         //                      .export
		.TD_RESET                 (video_in_TD_RESET),                            //                      .export
		.overflow_flag            (video_in_overflow_flag)                        //                      .export
	);

	nios_system_Video_In_Chroma_Resampler video_in_chroma_resampler (
		.clk                      (sys_clk),                                                      //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                               //    clock_reset_reset.reset
		.stream_in_startofpacket  (video_in_avalon_decoder_source_startofpacket),                 //   avalon_chroma_sink.startofpacket
		.stream_in_endofpacket    (video_in_avalon_decoder_source_endofpacket),                   //                     .endofpacket
		.stream_in_valid          (video_in_avalon_decoder_source_valid),                         //                     .valid
		.stream_in_ready          (video_in_avalon_decoder_source_ready),                         //                     .ready
		.stream_in_data           (video_in_avalon_decoder_source_data),                          //                     .data
		.stream_out_ready         (video_in_chroma_resampler_avalon_chroma_source_ready),         // avalon_chroma_source.ready
		.stream_out_startofpacket (video_in_chroma_resampler_avalon_chroma_source_startofpacket), //                     .startofpacket
		.stream_out_endofpacket   (video_in_chroma_resampler_avalon_chroma_source_endofpacket),   //                     .endofpacket
		.stream_out_valid         (video_in_chroma_resampler_avalon_chroma_source_valid),         //                     .valid
		.stream_out_data          (video_in_chroma_resampler_avalon_chroma_source_data)           //                     .data
	);

	nios_system_Video_In_CSC video_in_csc (
		.clk                      (sys_clk),                                                      //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                               // clock_reset_reset.reset
		.stream_in_startofpacket  (video_in_chroma_resampler_avalon_chroma_source_startofpacket), //   avalon_csc_sink.startofpacket
		.stream_in_endofpacket    (video_in_chroma_resampler_avalon_chroma_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (video_in_chroma_resampler_avalon_chroma_source_valid),         //                  .valid
		.stream_in_ready          (video_in_chroma_resampler_avalon_chroma_source_ready),         //                  .ready
		.stream_in_data           (video_in_chroma_resampler_avalon_chroma_source_data),          //                  .data
		.stream_out_ready         (video_in_csc_avalon_csc_source_ready),                         // avalon_csc_source.ready
		.stream_out_startofpacket (video_in_csc_avalon_csc_source_startofpacket),                 //                  .startofpacket
		.stream_out_endofpacket   (video_in_csc_avalon_csc_source_endofpacket),                   //                  .endofpacket
		.stream_out_valid         (video_in_csc_avalon_csc_source_valid),                         //                  .valid
		.stream_out_data          (video_in_csc_avalon_csc_source_data)                           //                  .data
	);

	nios_system_Video_In_RGB_Resampler video_in_rgb_resampler (
		.clk                      (sys_clk),                                                //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                         // clock_reset_reset.reset
		.stream_in_startofpacket  (video_in_csc_avalon_csc_source_startofpacket),           //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_in_csc_avalon_csc_source_endofpacket),             //                  .endofpacket
		.stream_in_valid          (video_in_csc_avalon_csc_source_valid),                   //                  .valid
		.stream_in_ready          (video_in_csc_avalon_csc_source_ready),                   //                  .ready
		.stream_in_data           (video_in_csc_avalon_csc_source_data),                    //                  .data
		.stream_out_ready         (video_in_rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (video_in_rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (video_in_rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (video_in_rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (video_in_rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	nios_system_Video_In_Clipper video_in_clipper (
		.clk                      (sys_clk),                                                //           clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                         //     clock_reset_reset.reset
		.stream_in_data           (video_in_rgb_resampler_avalon_rgb_source_data),          //   avalon_clipper_sink.data
		.stream_in_startofpacket  (video_in_rgb_resampler_avalon_rgb_source_startofpacket), //                      .startofpacket
		.stream_in_endofpacket    (video_in_rgb_resampler_avalon_rgb_source_endofpacket),   //                      .endofpacket
		.stream_in_valid          (video_in_rgb_resampler_avalon_rgb_source_valid),         //                      .valid
		.stream_in_ready          (video_in_rgb_resampler_avalon_rgb_source_ready),         //                      .ready
		.stream_out_ready         (video_in_clipper_avalon_clipper_source_ready),           // avalon_clipper_source.ready
		.stream_out_data          (video_in_clipper_avalon_clipper_source_data),            //                      .data
		.stream_out_startofpacket (video_in_clipper_avalon_clipper_source_startofpacket),   //                      .startofpacket
		.stream_out_endofpacket   (video_in_clipper_avalon_clipper_source_endofpacket),     //                      .endofpacket
		.stream_out_valid         (video_in_clipper_avalon_clipper_source_valid)            //                      .valid
	);

	nios_system_Video_In_Scaler video_in_scaler (
		.clk                      (sys_clk),                                              //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                       //    clock_reset_reset.reset
		.stream_in_startofpacket  (video_in_clipper_avalon_clipper_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_in_clipper_avalon_clipper_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_in_clipper_avalon_clipper_source_valid),         //                     .valid
		.stream_in_ready          (video_in_clipper_avalon_clipper_source_ready),         //                     .ready
		.stream_in_data           (video_in_clipper_avalon_clipper_source_data),          //                     .data
		.stream_out_ready         (video_in_scaler_avalon_scaler_source_ready),           // avalon_scaler_source.ready
		.stream_out_startofpacket (video_in_scaler_avalon_scaler_source_startofpacket),   //                     .startofpacket
		.stream_out_endofpacket   (video_in_scaler_avalon_scaler_source_endofpacket),     //                     .endofpacket
		.stream_out_valid         (video_in_scaler_avalon_scaler_source_valid),           //                     .valid
		.stream_out_data          (video_in_scaler_avalon_scaler_source_data)             //                     .data
	);

	nios_system_Camera_Config camera_config (
		.clk         (sys_clk),                                                                         //            clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                                  //      clock_reset_reset.reset
		.address     (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address),     // avalon_av_config_slave.address
		.byteenable  (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),  //                       .byteenable
		.read        (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read),        //                       .read
		.write       (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write),       //                       .write
		.writedata   (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),   //                       .writedata
		.readdata    (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),    //                       .readdata
		.waitrequest (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest), //                       .waitrequest
		.I2C_SDAT    (camera_config_I2C_SDAT),                                                          //     external_interface.export
		.I2C_SCLK    (camera_config_I2C_SCLK),                                                          //                       .export
		.exposure    (camera_config_exposure)                                                           //                       .export
	);

	nios_system_Camera_In camera_in (
		.clk                      (sys_clk),                                       //           clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                //     clock_reset_reset.reset
		.stream_out_ready         (camera_in_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (camera_in_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (camera_in_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (camera_in_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (camera_in_avalon_decoder_source_data),          //                      .data
		.PIXEL_CLK                (camera_in_PIXEL_CLK),                           //    external_interface.export
		.LINE_VALID               (camera_in_LINE_VALID),                          //                      .export
		.FRAME_VALID              (camera_in_FRAME_VALID),                         //                      .export
		.pixel_clk_reset          (camera_in_pixel_clk_reset),                     //                      .export
		.PIXEL_DATA               (camera_in_PIXEL_DATA)                           //                      .export
	);

	nios_system_Camera_Bayer_Resampler camera_bayer_resampler (
		.clk                      (sys_clk),                                                  //         clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                           //   clock_reset_reset.reset
		.stream_in_data           (camera_in_avalon_decoder_source_data),                     //   avalon_bayer_sink.data
		.stream_in_startofpacket  (camera_in_avalon_decoder_source_startofpacket),            //                    .startofpacket
		.stream_in_endofpacket    (camera_in_avalon_decoder_source_endofpacket),              //                    .endofpacket
		.stream_in_valid          (camera_in_avalon_decoder_source_valid),                    //                    .valid
		.stream_in_ready          (camera_in_avalon_decoder_source_ready),                    //                    .ready
		.stream_out_ready         (camera_bayer_resampler_avalon_bayer_source_ready),         // avalon_bayer_source.ready
		.stream_out_data          (camera_bayer_resampler_avalon_bayer_source_data),          //                    .data
		.stream_out_startofpacket (camera_bayer_resampler_avalon_bayer_source_startofpacket), //                    .startofpacket
		.stream_out_endofpacket   (camera_bayer_resampler_avalon_bayer_source_endofpacket),   //                    .endofpacket
		.stream_out_valid         (camera_bayer_resampler_avalon_bayer_source_valid)          //                    .valid
	);

	nios_system_Camera_Scaler camera_scaler (
		.clk                      (sys_clk),                                                  //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                           //    clock_reset_reset.reset
		.stream_in_startofpacket  (camera_bayer_resampler_avalon_bayer_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (camera_bayer_resampler_avalon_bayer_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (camera_bayer_resampler_avalon_bayer_source_valid),         //                     .valid
		.stream_in_ready          (camera_bayer_resampler_avalon_bayer_source_ready),         //                     .ready
		.stream_in_data           (camera_bayer_resampler_avalon_bayer_source_data),          //                     .data
		.stream_out_ready         (camera_scaler_avalon_scaler_source_ready),                 // avalon_scaler_source.ready
		.stream_out_startofpacket (camera_scaler_avalon_scaler_source_startofpacket),         //                     .startofpacket
		.stream_out_endofpacket   (camera_scaler_avalon_scaler_source_endofpacket),           //                     .endofpacket
		.stream_out_valid         (camera_scaler_avalon_scaler_source_valid),                 //                     .valid
		.stream_out_data          (camera_scaler_avalon_scaler_source_data)                   //                     .data
	);

	nios_system_Camera_Clipper camera_clipper (
		.clk                      (sys_clk),                                            //           clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                     //     clock_reset_reset.reset
		.stream_in_data           (camera_scaler_avalon_scaler_source_data),            //   avalon_clipper_sink.data
		.stream_in_startofpacket  (camera_scaler_avalon_scaler_source_startofpacket),   //                      .startofpacket
		.stream_in_endofpacket    (camera_scaler_avalon_scaler_source_endofpacket),     //                      .endofpacket
		.stream_in_valid          (camera_scaler_avalon_scaler_source_valid),           //                      .valid
		.stream_in_ready          (camera_scaler_avalon_scaler_source_ready),           //                      .ready
		.stream_out_ready         (camera_clipper_avalon_clipper_source_ready),         // avalon_clipper_source.ready
		.stream_out_data          (camera_clipper_avalon_clipper_source_data),          //                      .data
		.stream_out_startofpacket (camera_clipper_avalon_clipper_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (camera_clipper_avalon_clipper_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (camera_clipper_avalon_clipper_source_valid)          //                      .valid
	);

	nios_system_Video_In_RGB_Resampler camera_rgb_resampler (
		.clk                      (sys_clk),                                              //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                       // clock_reset_reset.reset
		.stream_in_startofpacket  (camera_clipper_avalon_clipper_source_startofpacket),   //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (camera_clipper_avalon_clipper_source_endofpacket),     //                  .endofpacket
		.stream_in_valid          (camera_clipper_avalon_clipper_source_valid),           //                  .valid
		.stream_in_ready          (camera_clipper_avalon_clipper_source_ready),           //                  .ready
		.stream_in_data           (camera_clipper_avalon_clipper_source_data),            //                  .data
		.stream_out_ready         (camera_rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (camera_rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (camera_rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (camera_rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (camera_rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	nios_system_LCD_Controller lcd_controller (
		.clk           (external_clocks_vga_clk_33_clk),                            //        clock_reset.clk
		.reset         (rst_controller_004_reset_out_reset),                        //  clock_reset_reset.reset
		.data          (lcd_dual_clock_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (lcd_dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (lcd_dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (lcd_dual_clock_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (lcd_dual_clock_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (lcd_controller_external_interface_CLK),                     // external_interface.export
		.VGA_HS        (lcd_controller_external_interface_HS),                      //                   .export
		.VGA_VS        (lcd_controller_external_interface_VS),                      //                   .export
		.VGA_DATA_EN   (lcd_controller_external_interface_DATA_EN),                 //                   .export
		.VGA_R         (lcd_controller_external_interface_R),                       //                   .export
		.VGA_G         (lcd_controller_external_interface_G),                       //                   .export
		.VGA_B         (lcd_controller_external_interface_B)                        //                   .export
	);

	nios_system_LCD_RGB_Resampler lcd_rgb_resampler (
		.clk                      (sys_clk),                                              //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                       // clock_reset_reset.reset
		.stream_in_startofpacket  (lcd_dma_controller_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (lcd_dma_controller_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (lcd_dma_controller_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (lcd_dma_controller_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (lcd_dma_controller_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (lcd_rgb_resampler_avalon_rgb_source_ready),            // avalon_rgb_source.ready
		.stream_out_startofpacket (lcd_rgb_resampler_avalon_rgb_source_startofpacket),    //                  .startofpacket
		.stream_out_endofpacket   (lcd_rgb_resampler_avalon_rgb_source_endofpacket),      //                  .endofpacket
		.stream_out_valid         (lcd_rgb_resampler_avalon_rgb_source_valid),            //                  .valid
		.stream_out_data          (lcd_rgb_resampler_avalon_rgb_source_data)              //                  .data
	);

	nios_system_LCD_Scalar lcd_scalar (
		.clk                      (sys_clk),                                           //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                    //    clock_reset_reset.reset
		.stream_in_startofpacket  (lcd_rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (lcd_rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (lcd_rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (lcd_rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (lcd_rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (lcd_scalar_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (lcd_scalar_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (lcd_scalar_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (lcd_scalar_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (lcd_scalar_avalon_scaler_source_data)               //                     .data
	);

	nios_system_LCD_Dual_Clock_FIFO lcd_dual_clock_fifo (
		.clk_stream_in            (sys_clk),                                                   //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                            //   clock_stream_in_reset.reset
		.clk_stream_out           (external_clocks_vga_clk_33_clk),                            //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_004_reset_out_reset),                        //  clock_stream_out_reset.reset
		.stream_in_ready          (lcd_alpha_blender_avalon_blended_source_ready),             //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (lcd_alpha_blender_avalon_blended_source_startofpacket),     //                        .startofpacket
		.stream_in_endofpacket    (lcd_alpha_blender_avalon_blended_source_endofpacket),       //                        .endofpacket
		.stream_in_valid          (lcd_alpha_blender_avalon_blended_source_valid),             //                        .valid
		.stream_in_data           (lcd_alpha_blender_avalon_blended_source_data),              //                        .data
		.stream_out_ready         (lcd_dual_clock_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (lcd_dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (lcd_dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (lcd_dual_clock_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (lcd_dual_clock_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	nios_system_Video_In_DMA_Controller video_in_dma_controller (
		.clk                  (sys_clk),                                                                                    //              clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                             //        clock_reset_reset.reset
		.stream_data          (video_in_scaler_avalon_scaler_source_data),                                                  //          avalon_dma_sink.data
		.stream_startofpacket (video_in_scaler_avalon_scaler_source_startofpacket),                                         //                         .startofpacket
		.stream_endofpacket   (video_in_scaler_avalon_scaler_source_endofpacket),                                           //                         .endofpacket
		.stream_valid         (video_in_scaler_avalon_scaler_source_valid),                                                 //                         .valid
		.stream_ready         (video_in_scaler_avalon_scaler_source_ready),                                                 //                         .ready
		.slave_address        (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable), //                         .byteenable
		.slave_read           (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),       //                         .read
		.slave_write          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),      //                         .write
		.slave_writedata      (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),  //                         .writedata
		.slave_readdata       (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),   //                         .readdata
		.master_address       (video_in_dma_controller_avalon_dma_master_address),                                          //        avalon_dma_master.address
		.master_waitrequest   (video_in_dma_controller_avalon_dma_master_waitrequest),                                      //                         .waitrequest
		.master_write         (video_in_dma_controller_avalon_dma_master_write),                                            //                         .write
		.master_writedata     (video_in_dma_controller_avalon_dma_master_writedata)                                         //                         .writedata
	);

	nios_system_Camera_DMA_Controller camera_dma_controller (
		.clk                  (sys_clk),                                                                                  //              clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                           //        clock_reset_reset.reset
		.stream_data          (camera_rgb_resampler_avalon_rgb_source_data),                                              //          avalon_dma_sink.data
		.stream_startofpacket (camera_rgb_resampler_avalon_rgb_source_startofpacket),                                     //                         .startofpacket
		.stream_endofpacket   (camera_rgb_resampler_avalon_rgb_source_endofpacket),                                       //                         .endofpacket
		.stream_valid         (camera_rgb_resampler_avalon_rgb_source_valid),                                             //                         .valid
		.stream_ready         (camera_rgb_resampler_avalon_rgb_source_ready),                                             //                         .ready
		.slave_address        (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable), //                         .byteenable
		.slave_read           (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),       //                         .read
		.slave_write          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),      //                         .write
		.slave_writedata      (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),  //                         .writedata
		.slave_readdata       (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),   //                         .readdata
		.master_address       (camera_dma_controller_avalon_dma_master_address),                                          //        avalon_dma_master.address
		.master_waitrequest   (camera_dma_controller_avalon_dma_master_waitrequest),                                      //                         .waitrequest
		.master_write         (camera_dma_controller_avalon_dma_master_write),                                            //                         .write
		.master_writedata     (camera_dma_controller_avalon_dma_master_writedata)                                         //                         .writedata
	);

	nios_system_Accelerometer accelerometer (
		.clk           (sys_clk),                                                                                      //                         clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                                               //                   clock_reset_reset.reset
		.address       (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_address),     // avalon_accelerometer_spi_mode_slave.address
		.byteenable    (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_byteenable),  //                                    .byteenable
		.read          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_read),        //                                    .read
		.write         (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_write),       //                                    .write
		.writedata     (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_writedata),   //                                    .writedata
		.readdata      (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_readdata),    //                                    .readdata
		.waitrequest   (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_waitrequest), //                                    .waitrequest
		.irq           (irq_mapper_receiver9_irq),                                                                     //                           interrupt.irq
		.I2C_SDAT      (accelerometer_I2C_SDAT),                                                                       //                  external_interface.export
		.I2C_SCLK      (accelerometer_I2C_SCLK),                                                                       //                                    .export
		.G_SENSOR_CS_N (accelerometer_G_SENSOR_CS_N),                                                                  //                                    .export
		.G_SENSOR_INT  (accelerometer_G_SENSOR_INT)                                                                    //                                    .export
	);

	nios_system_USB usb (
		.clk        (sys_clk),                                                        //        clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                 //  clock_reset_reset.reset
		.address    (usb_avalon_usb_slave_translator_avalon_anti_slave_0_address),    //   avalon_usb_slave.address
		.chipselect (usb_avalon_usb_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.read       (usb_avalon_usb_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write      (usb_avalon_usb_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata  (usb_avalon_usb_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata   (usb_avalon_usb_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver10_irq),                                      //          interrupt.irq
		.OTG_INT1   (usb_INT1),                                                       // external_interface.export
		.OTG_DATA   (usb_DATA),                                                       //                   .export
		.OTG_RST_N  (usb_RST_N),                                                      //                   .export
		.OTG_ADDR   (usb_ADDR),                                                       //                   .export
		.OTG_CS_N   (usb_CS_N),                                                       //                   .export
		.OTG_RD_N   (usb_RD_N),                                                       //                   .export
		.OTG_WR_N   (usb_WR_N),                                                       //                   .export
		.OTG_INT0   (usb_INT0)                                                        //                   .export
	);

	nios_system_LCD_Char_Buffer lcd_char_buffer (
		.clk                  (sys_clk),                                                                             //               clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                      //         clock_reset_reset.reset
		.ctrl_address         (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable), //                          .byteenable
		.ctrl_chipselect      (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect), //                          .chipselect
		.ctrl_read            (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read),       //                          .read
		.ctrl_write           (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write),      //                          .write
		.ctrl_writedata       (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),  //                          .writedata
		.ctrl_readdata        (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),   //                          .readdata
		.buf_byteenable       (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),  //                          .chipselect
		.buf_read             (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),        //                          .read
		.buf_write            (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),       //                          .write
		.buf_writedata        (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.buf_readdata         (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.buf_waitrequest      (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.buf_address          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),     //                          .address
		.stream_ready         (lcd_char_buffer_avalon_char_source_ready),                                            //        avalon_char_source.ready
		.stream_startofpacket (lcd_char_buffer_avalon_char_source_startofpacket),                                    //                          .startofpacket
		.stream_endofpacket   (lcd_char_buffer_avalon_char_source_endofpacket),                                      //                          .endofpacket
		.stream_valid         (lcd_char_buffer_avalon_char_source_valid),                                            //                          .valid
		.stream_data          (lcd_char_buffer_avalon_char_source_data)                                              //                          .data
	);

	nios_system_VGA_Alpha_Blender lcd_alpha_blender (
		.clk                      (sys_clk),                                               //            clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                        //      clock_reset_reset.reset
		.foreground_data          (lcd_char_buffer_avalon_char_source_data),               // avalon_foreground_sink.data
		.foreground_startofpacket (lcd_char_buffer_avalon_char_source_startofpacket),      //                       .startofpacket
		.foreground_endofpacket   (lcd_char_buffer_avalon_char_source_endofpacket),        //                       .endofpacket
		.foreground_valid         (lcd_char_buffer_avalon_char_source_valid),              //                       .valid
		.foreground_ready         (lcd_char_buffer_avalon_char_source_ready),              //                       .ready
		.background_data          (lcd_scalar_avalon_scaler_source_data),                  // avalon_background_sink.data
		.background_startofpacket (lcd_scalar_avalon_scaler_source_startofpacket),         //                       .startofpacket
		.background_endofpacket   (lcd_scalar_avalon_scaler_source_endofpacket),           //                       .endofpacket
		.background_valid         (lcd_scalar_avalon_scaler_source_valid),                 //                       .valid
		.background_ready         (lcd_scalar_avalon_scaler_source_ready),                 //                       .ready
		.output_ready             (lcd_alpha_blender_avalon_blended_source_ready),         //  avalon_blended_source.ready
		.output_data              (lcd_alpha_blender_avalon_blended_source_data),          //                       .data
		.output_startofpacket     (lcd_alpha_blender_avalon_blended_source_startofpacket), //                       .startofpacket
		.output_endofpacket       (lcd_alpha_blender_avalon_blended_source_endofpacket),   //                       .endofpacket
		.output_valid             (lcd_alpha_blender_avalon_blended_source_valid)          //                       .valid
	);

	nios_system_enet enet (
		.clk           (sys_clk),                                                      // control_port_clock_connection.clk
		.reset         (rst_controller_005_reset_out_reset),                           //              reset_connection.reset
		.address       (enet_control_port_translator_avalon_anti_slave_0_address),     //                  control_port.address
		.readdata      (enet_control_port_translator_avalon_anti_slave_0_readdata),    //                              .readdata
		.read          (enet_control_port_translator_avalon_anti_slave_0_read),        //                              .read
		.writedata     (enet_control_port_translator_avalon_anti_slave_0_writedata),   //                              .writedata
		.write         (enet_control_port_translator_avalon_anti_slave_0_write),       //                              .write
		.waitrequest   (enet_control_port_translator_avalon_anti_slave_0_waitrequest), //                              .waitrequest
		.tx_clk        (enet_pcs_mac_tx_clk),                                          //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (enet_pcs_mac_rx_clk),                                          //   pcs_mac_rx_clock_connection.clk
		.set_10        (enet_mac_status_set_10),                                       //         mac_status_connection.set_10
		.set_1000      (enet_mac_status_set_1000),                                     //                              .set_1000
		.eth_mode      (enet_mac_status_eth_mode),                                     //                              .eth_mode
		.ena_10        (enet_mac_status_ena_10),                                       //                              .ena_10
		.rgmii_in      (enet_mac_rgmii_rgmii_in),                                      //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (enet_mac_rgmii_rgmii_out),                                     //                              .rgmii_out
		.rx_control    (enet_mac_rgmii_rx_control),                                    //                              .rx_control
		.tx_control    (enet_mac_rgmii_tx_control),                                    //                              .tx_control
		.ff_rx_clk     (sys_clk),                                                      //     transmit_clock_connection.clk
		.ff_tx_clk     (sys_clk),                                                      //      receive_clock_connection.clk
		.ff_rx_data    (enet_receive_data),                                            //                       receive.data
		.ff_rx_eop     (enet_receive_endofpacket),                                     //                              .endofpacket
		.rx_err        (enet_receive_error),                                           //                              .error
		.ff_rx_mod     (enet_receive_empty),                                           //                              .empty
		.ff_rx_rdy     (enet_receive_ready),                                           //                              .ready
		.ff_rx_sop     (enet_receive_startofpacket),                                   //                              .startofpacket
		.ff_rx_dval    (enet_receive_valid),                                           //                              .valid
		.ff_tx_data    (avalon_st_adapter_001_out_0_data),                             //                      transmit.data
		.ff_tx_eop     (avalon_st_adapter_001_out_0_endofpacket),                      //                              .endofpacket
		.ff_tx_err     (avalon_st_adapter_001_out_0_error),                            //                              .error
		.ff_tx_mod     (avalon_st_adapter_001_out_0_empty),                            //                              .empty
		.ff_tx_rdy     (avalon_st_adapter_001_out_0_ready),                            //                              .ready
		.ff_tx_sop     (avalon_st_adapter_001_out_0_startofpacket),                    //                              .startofpacket
		.ff_tx_wren    (avalon_st_adapter_001_out_0_valid),                            //                              .valid
		.mdc           (enet_mac_mdio_mdc),                                            //           mac_mdio_connection.mdc
		.mdio_in       (enet_mac_mdio_mdio_in),                                        //                              .mdio_in
		.mdio_out      (enet_mac_mdio_mdio_out),                                       //                              .mdio_out
		.mdio_oen      (enet_mac_mdio_mdio_oen),                                       //                              .mdio_oen
		.xon_gen       (enet_mac_misc_xon_gen),                                        //           mac_misc_connection.xon_gen
		.xoff_gen      (enet_mac_misc_xoff_gen),                                       //                              .xoff_gen
		.magic_wakeup  (enet_mac_misc_magic_wakeup),                                   //                              .magic_wakeup
		.magic_sleep_n (enet_mac_misc_magic_sleep_n),                                  //                              .magic_sleep_n
		.ff_tx_crc_fwd (enet_mac_misc_ff_tx_crc_fwd),                                  //                              .ff_tx_crc_fwd
		.ff_tx_septy   (enet_mac_misc_ff_tx_septy),                                    //                              .ff_tx_septy
		.tx_ff_uflow   (enet_mac_misc_tx_ff_uflow),                                    //                              .tx_ff_uflow
		.ff_tx_a_full  (enet_mac_misc_ff_tx_a_full),                                   //                              .ff_tx_a_full
		.ff_tx_a_empty (enet_mac_misc_ff_tx_a_empty),                                  //                              .ff_tx_a_empty
		.rx_err_stat   (enet_mac_misc_rx_err_stat),                                    //                              .rx_err_stat
		.rx_frm_type   (enet_mac_misc_rx_frm_type),                                    //                              .rx_frm_type
		.ff_rx_dsav    (enet_mac_misc_ff_rx_dsav),                                     //                              .ff_rx_dsav
		.ff_rx_a_full  (enet_mac_misc_ff_rx_a_full),                                   //                              .ff_rx_a_full
		.ff_rx_a_empty (enet_mac_misc_ff_rx_a_empty)                                   //                              .ff_rx_a_empty
	);

	nios_system_descriptor_memory descriptor_memory (
		.clk        (sys_clk),                                                        //   clk1.clk
		.address    (descriptor_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (descriptor_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_005_reset_out_reset),                             // reset1.reset
		.reset_req  (rst_controller_005_reset_out_reset_req)                          //       .reset_req
	);

	nios_system_packet_memory packet_memory (
		.clk        (sys_clk),                                                    //   clk1.clk
		.address    (packet_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (packet_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (packet_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (packet_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (packet_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (packet_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (packet_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_005_reset_out_reset),                         // reset1.reset
		.reset_req  (rst_controller_005_reset_out_reset_req)                      //       .reset_req
	);

	nios_system_LCD_DMA_Controller lcd_dma_controller (
		.clk                  (sys_clk),                                                                               //              clock_reset.clk
		.reset                (cpu_jtag_debug_module_reset_reset),                                                     //        clock_reset_reset.reset
		.master_address       (lcd_dma_controller_avalon_dma_master_address),                                          //        avalon_dma_master.address
		.master_waitrequest   (lcd_dma_controller_avalon_dma_master_waitrequest),                                      //                         .waitrequest
		.master_arbiterlock   (lcd_dma_controller_avalon_dma_master_lock),                                             //                         .lock
		.master_read          (lcd_dma_controller_avalon_dma_master_read),                                             //                         .read
		.master_readdata      (lcd_dma_controller_avalon_dma_master_readdata),                                         //                         .readdata
		.master_readdatavalid (lcd_dma_controller_avalon_dma_master_readdatavalid),                                    //                         .readdatavalid
		.slave_address        (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable), //                         .byteenable
		.slave_read           (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),       //                         .read
		.slave_write          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),      //                         .write
		.slave_writedata      (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),  //                         .writedata
		.slave_readdata       (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),   //                         .readdata
		.stream_ready         (lcd_dma_controller_avalon_pixel_source_ready),                                          //      avalon_pixel_source.ready
		.stream_data          (lcd_dma_controller_avalon_pixel_source_data),                                           //                         .data
		.stream_startofpacket (lcd_dma_controller_avalon_pixel_source_startofpacket),                                  //                         .startofpacket
		.stream_endofpacket   (lcd_dma_controller_avalon_pixel_source_endofpacket),                                    //                         .endofpacket
		.stream_valid         (lcd_dma_controller_avalon_pixel_source_valid)                                           //                         .valid
	);

	nios_system_VGA_DMA_Controller vga_dma_controller (
		.clk                  (sys_clk),                                                                               //              clock_reset.clk
		.reset                (cpu_jtag_debug_module_reset_reset),                                                     //        clock_reset_reset.reset
		.master_address       (vga_dma_controller_avalon_dma_master_address),                                          //        avalon_dma_master.address
		.master_waitrequest   (vga_dma_controller_avalon_dma_master_waitrequest),                                      //                         .waitrequest
		.master_arbiterlock   (vga_dma_controller_avalon_dma_master_lock),                                             //                         .lock
		.master_read          (vga_dma_controller_avalon_dma_master_read),                                             //                         .read
		.master_readdata      (vga_dma_controller_avalon_dma_master_readdata),                                         //                         .readdata
		.master_readdatavalid (vga_dma_controller_avalon_dma_master_readdatavalid),                                    //                         .readdatavalid
		.slave_address        (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable), //                         .byteenable
		.slave_read           (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),       //                         .read
		.slave_write          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),      //                         .write
		.slave_writedata      (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),  //                         .writedata
		.slave_readdata       (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),   //                         .readdata
		.stream_ready         (vga_dma_controller_avalon_pixel_source_ready),                                          //      avalon_pixel_source.ready
		.stream_data          (vga_dma_controller_avalon_pixel_source_data),                                           //                         .data
		.stream_startofpacket (vga_dma_controller_avalon_pixel_source_startofpacket),                                  //                         .startofpacket
		.stream_endofpacket   (vga_dma_controller_avalon_pixel_source_endofpacket),                                    //                         .endofpacket
		.stream_valid         (vga_dma_controller_avalon_pixel_source_valid)                                           //                         .valid
	);

	VideoConferencing_DMA videoconferencing_dma_0 (
		.slave_chipselect   (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_chipselect), //            avalon_slave.chipselect
		.slave_writedata    (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_writedata),  //                        .writedata
		.slave_readdata     (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_readdata),   //                        .readdata
		.slave_read         (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_read),       //                        .read
		.slave_address      (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_address),    //                        .address
		.slave_write        (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_write),      //                        .write
		.master_waitrequest (videoconferencing_dma_0_avalon_master_waitrequest),                              //           avalon_master.waitrequest
		.master_address     (videoconferencing_dma_0_avalon_master_address),                                  //                        .address
		.master_write       (videoconferencing_dma_0_avalon_master_write),                                    //                        .write
		.master_byteenable  (videoconferencing_dma_0_avalon_master_byteenable),                               //                        .byteenable
		.master_writedata   (videoconferencing_dma_0_avalon_master_writedata),                                //                        .writedata
		.LEDR_conduit       (videoconferencing_dma_conduit_LEDR_conduit),                                     //             conduit_end.export
		.LEDG_conduit       (videoconferencing_dma_conduit_LEDG_conduit),                                     //                        .export
		.HEX0_conduit       (videoconferencing_dma_conduit_HEX0_conduit),                                     //                        .export
		.HEX1_conduit       (videoconferencing_dma_conduit_HEX1_conduit),                                     //                        .export
		.HEX2_conduit       (videoconferencing_dma_conduit_HEX2_conduit),                                     //                        .export
		.HEX3_conduit       (videoconferencing_dma_conduit_HEX3_conduit),                                     //                        .export
		.HEX4_conduit       (videoconferencing_dma_conduit_HEX4_conduit),                                     //                        .export
		.HEX5_conduit       (videoconferencing_dma_conduit_HEX5_conduit),                                     //                        .export
		.HEX6_conduit       (videoconferencing_dma_conduit_HEX6_conduit),                                     //                        .export
		.HEX7_conduit       (videoconferencing_dma_conduit_HEX7_conduit),                                     //                        .export
		.SW_conduit         (videoconferencing_dma_conduit_SW_conduit),                                       //                        .export
		.clk                (sys_clk),                                                                        //              clock_sink.clk
		.eth_rx_mod         (avalon_st_adapter_out_0_channel),                                                //   avalon_streaming_sink.channel
		.eth_rx_data        (avalon_st_adapter_out_0_data),                                                   //                        .data
		.eth_rx_sop         (avalon_st_adapter_out_0_startofpacket),                                          //                        .startofpacket
		.eth_rx_error       (avalon_st_adapter_out_0_error),                                                  //                        .error
		.eth_rx_dval        (avalon_st_adapter_out_0_valid),                                                  //                        .valid
		.eth_rx_rdy         (avalon_st_adapter_out_0_ready),                                                  //                        .ready
		.eth_rx_eop         (avalon_st_adapter_out_0_endofpacket),                                            //                        .endofpacket
		.eth_tx_error       (videoconferencing_dma_0_avalon_streaming_source_error),                          // avalon_streaming_source.error
		.eth_tx_rdy         (videoconferencing_dma_0_avalon_streaming_source_ready),                          //                        .ready
		.eth_tx_data        (videoconferencing_dma_0_avalon_streaming_source_data),                           //                        .data
		.eth_tx_mod         (videoconferencing_dma_0_avalon_streaming_source_channel),                        //                        .channel
		.eth_tx_wren        (videoconferencing_dma_0_avalon_streaming_source_valid),                          //                        .valid
		.eth_tx_sop         (videoconferencing_dma_0_avalon_streaming_source_startofpacket),                  //                        .startofpacket
		.eth_tx_eop         (videoconferencing_dma_0_avalon_streaming_source_endofpacket),                    //                        .endofpacket
		.resetn             (~rst_controller_006_reset_out_reset)                                             //              reset_sink.reset_n
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) cpu_custom_instruction_master_translator (
		.ci_slave_result         (),                                                                 //        ci_slave.result
		.ci_slave_multi_clk      (cpu_custom_instruction_master_clk),                                //                .clk
		.ci_slave_multi_reset    (cpu_custom_instruction_master_reset),                              //                .reset
		.ci_slave_multi_clken    (cpu_custom_instruction_master_clk_en),                             //                .clk_en
		.ci_slave_multi_start    (cpu_custom_instruction_master_start),                              //                .start
		.ci_slave_multi_done     (cpu_custom_instruction_master_done),                               //                .done
		.ci_slave_multi_dataa    (cpu_custom_instruction_master_multi_dataa),                        //                .multi_dataa
		.ci_slave_multi_datab    (cpu_custom_instruction_master_multi_datab),                        //                .multi_datab
		.ci_slave_multi_result   (cpu_custom_instruction_master_multi_result),                       //                .multi_result
		.ci_slave_multi_n        (cpu_custom_instruction_master_multi_n),                            //                .multi_n
		.ci_slave_multi_readra   (cpu_custom_instruction_master_multi_readra),                       //                .multi_readra
		.ci_slave_multi_readrb   (cpu_custom_instruction_master_multi_readrb),                       //                .multi_readrb
		.ci_slave_multi_writerc  (cpu_custom_instruction_master_multi_writerc),                      //                .multi_writerc
		.ci_slave_multi_a        (cpu_custom_instruction_master_multi_a),                            //                .multi_a
		.ci_slave_multi_b        (cpu_custom_instruction_master_multi_b),                            //                .multi_b
		.ci_slave_multi_c        (cpu_custom_instruction_master_multi_c),                            //                .multi_c
		.comb_ci_master_result   (),                                                                 //  comb_ci_master.result
		.multi_ci_master_clk     (cpu_custom_instruction_master_translator_multi_ci_master_clk),     // multi_ci_master.clk
		.multi_ci_master_reset   (cpu_custom_instruction_master_translator_multi_ci_master_reset),   //                .reset
		.multi_ci_master_clken   (cpu_custom_instruction_master_translator_multi_ci_master_clk_en),  //                .clk_en
		.multi_ci_master_start   (cpu_custom_instruction_master_translator_multi_ci_master_start),   //                .start
		.multi_ci_master_done    (cpu_custom_instruction_master_translator_multi_ci_master_done),    //                .done
		.multi_ci_master_dataa   (cpu_custom_instruction_master_translator_multi_ci_master_dataa),   //                .dataa
		.multi_ci_master_datab   (cpu_custom_instruction_master_translator_multi_ci_master_datab),   //                .datab
		.multi_ci_master_result  (cpu_custom_instruction_master_translator_multi_ci_master_result),  //                .result
		.multi_ci_master_n       (cpu_custom_instruction_master_translator_multi_ci_master_n),       //                .n
		.multi_ci_master_readra  (cpu_custom_instruction_master_translator_multi_ci_master_readra),  //                .readra
		.multi_ci_master_readrb  (cpu_custom_instruction_master_translator_multi_ci_master_readrb),  //                .readrb
		.multi_ci_master_writerc (cpu_custom_instruction_master_translator_multi_ci_master_writerc), //                .writerc
		.multi_ci_master_a       (cpu_custom_instruction_master_translator_multi_ci_master_a),       //                .a
		.multi_ci_master_b       (cpu_custom_instruction_master_translator_multi_ci_master_b),       //                .b
		.multi_ci_master_c       (cpu_custom_instruction_master_translator_multi_ci_master_c),       //                .c
		.ci_slave_dataa          (32'b00000000000000000000000000000000),                             //     (terminated)
		.ci_slave_datab          (32'b00000000000000000000000000000000),                             //     (terminated)
		.ci_slave_n              (8'b00000000),                                                      //     (terminated)
		.ci_slave_readra         (1'b0),                                                             //     (terminated)
		.ci_slave_readrb         (1'b0),                                                             //     (terminated)
		.ci_slave_writerc        (1'b0),                                                             //     (terminated)
		.ci_slave_a              (5'b00000),                                                         //     (terminated)
		.ci_slave_b              (5'b00000),                                                         //     (terminated)
		.ci_slave_c              (5'b00000),                                                         //     (terminated)
		.ci_slave_ipending       (32'b00000000000000000000000000000000),                             //     (terminated)
		.ci_slave_estatus        (1'b0),                                                             //     (terminated)
		.comb_ci_master_dataa    (),                                                                 //     (terminated)
		.comb_ci_master_datab    (),                                                                 //     (terminated)
		.comb_ci_master_n        (),                                                                 //     (terminated)
		.comb_ci_master_readra   (),                                                                 //     (terminated)
		.comb_ci_master_readrb   (),                                                                 //     (terminated)
		.comb_ci_master_writerc  (),                                                                 //     (terminated)
		.comb_ci_master_a        (),                                                                 //     (terminated)
		.comb_ci_master_b        (),                                                                 //     (terminated)
		.comb_ci_master_c        (),                                                                 //     (terminated)
		.comb_ci_master_ipending (),                                                                 //     (terminated)
		.comb_ci_master_estatus  ()                                                                  //     (terminated)
	);

	nios_system_CPU_custom_instruction_master_multi_xconnect cpu_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa      (cpu_custom_instruction_master_translator_multi_ci_master_dataa),   //   ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_translator_multi_ci_master_datab),   //           .datab
		.ci_slave_result     (cpu_custom_instruction_master_translator_multi_ci_master_result),  //           .result
		.ci_slave_n          (cpu_custom_instruction_master_translator_multi_ci_master_n),       //           .n
		.ci_slave_readra     (cpu_custom_instruction_master_translator_multi_ci_master_readra),  //           .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_translator_multi_ci_master_readrb),  //           .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_translator_multi_ci_master_writerc), //           .writerc
		.ci_slave_a          (cpu_custom_instruction_master_translator_multi_ci_master_a),       //           .a
		.ci_slave_b          (cpu_custom_instruction_master_translator_multi_ci_master_b),       //           .b
		.ci_slave_c          (cpu_custom_instruction_master_translator_multi_ci_master_c),       //           .c
		.ci_slave_ipending   (),                                                                 //           .ipending
		.ci_slave_estatus    (),                                                                 //           .estatus
		.ci_slave_clk        (cpu_custom_instruction_master_translator_multi_ci_master_clk),     //           .clk
		.ci_slave_reset      (cpu_custom_instruction_master_translator_multi_ci_master_reset),   //           .reset
		.ci_slave_clken      (cpu_custom_instruction_master_translator_multi_ci_master_clk_en),  //           .clk_en
		.ci_slave_start      (cpu_custom_instruction_master_translator_multi_ci_master_start),   //           .start
		.ci_slave_done       (cpu_custom_instruction_master_translator_multi_ci_master_done),    //           .done
		.ci_master0_dataa    (cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa),    // ci_master0.dataa
		.ci_master0_datab    (cpu_custom_instruction_master_multi_xconnect_ci_master0_datab),    //           .datab
		.ci_master0_result   (cpu_custom_instruction_master_multi_xconnect_ci_master0_result),   //           .result
		.ci_master0_n        (cpu_custom_instruction_master_multi_xconnect_ci_master0_n),        //           .n
		.ci_master0_readra   (cpu_custom_instruction_master_multi_xconnect_ci_master0_readra),   //           .readra
		.ci_master0_readrb   (cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb),   //           .readrb
		.ci_master0_writerc  (cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc),  //           .writerc
		.ci_master0_a        (cpu_custom_instruction_master_multi_xconnect_ci_master0_a),        //           .a
		.ci_master0_b        (cpu_custom_instruction_master_multi_xconnect_ci_master0_b),        //           .b
		.ci_master0_c        (cpu_custom_instruction_master_multi_xconnect_ci_master0_c),        //           .c
		.ci_master0_ipending (cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending), //           .ipending
		.ci_master0_estatus  (cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus),  //           .estatus
		.ci_master0_clk      (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk),      //           .clk
		.ci_master0_reset    (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset),    //           .reset
		.ci_master0_clken    (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en),   //           .clk_en
		.ci_master0_start    (cpu_custom_instruction_master_multi_xconnect_ci_master0_start),    //           .start
		.ci_master0_done     (cpu_custom_instruction_master_multi_xconnect_ci_master0_done)      //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (2),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) cpu_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa     (cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab     (cpu_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result    (cpu_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n         (cpu_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra    (cpu_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb    (cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc   (cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a         (cpu_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b         (cpu_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c         (cpu_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending  (cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus   (cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk       (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken     (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset     (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start     (cpu_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done      (cpu_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result   (cpu_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n        (cpu_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk      (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra   (),                                                                       // (terminated)
		.ci_master_readrb   (),                                                                       // (terminated)
		.ci_master_writerc  (),                                                                       // (terminated)
		.ci_master_a        (),                                                                       // (terminated)
		.ci_master_b        (),                                                                       // (terminated)
		.ci_master_c        (),                                                                       // (terminated)
		.ci_master_ipending (),                                                                       // (terminated)
		.ci_master_estatus  ()                                                                        // (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                      (sys_clk),                                                                   //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (cpu_instruction_master_read),                                               //                          .read
		.av_readdata              (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_byteenable            (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_write                 (1'b0),                                                                      //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (29),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                      (sys_clk),                                                            //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address              (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_data_master_read),                                               //                          .read
		.av_readdata              (cpu_data_master_readdata),                                           //                          .readdata
		.av_write                 (cpu_data_master_write),                                              //                          .write
		.av_writedata             (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                               //               (terminated)
		.av_readdatavalid         (),                                                                   //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) video_in_dma_controller_avalon_dma_master_translator (
		.clk                      (sys_clk),                                                                                      //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                               //                     reset.reset
		.uav_address              (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (video_in_dma_controller_avalon_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (video_in_dma_controller_avalon_dma_master_waitrequest),                                        //                          .waitrequest
		.av_write                 (video_in_dma_controller_avalon_dma_master_write),                                              //                          .write
		.av_writedata             (video_in_dma_controller_avalon_dma_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                                         //               (terminated)
		.av_byteenable            (2'b11),                                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                         //               (terminated)
		.av_begintransfer         (1'b0),                                                                                         //               (terminated)
		.av_chipselect            (1'b0),                                                                                         //               (terminated)
		.av_read                  (1'b0),                                                                                         //               (terminated)
		.av_readdata              (),                                                                                             //               (terminated)
		.av_readdatavalid         (),                                                                                             //               (terminated)
		.av_lock                  (1'b0),                                                                                         //               (terminated)
		.av_debugaccess           (1'b0),                                                                                         //               (terminated)
		.uav_clken                (),                                                                                             //               (terminated)
		.av_clken                 (1'b1),                                                                                         //               (terminated)
		.uav_response             (2'b00),                                                                                        //               (terminated)
		.av_response              (),                                                                                             //               (terminated)
		.uav_writeresponserequest (),                                                                                             //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                         //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                         //               (terminated)
		.av_writeresponsevalid    ()                                                                                              //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) camera_dma_controller_avalon_dma_master_translator (
		.clk                      (sys_clk),                                                                                    //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                             //                     reset.reset
		.uav_address              (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (camera_dma_controller_avalon_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (camera_dma_controller_avalon_dma_master_waitrequest),                                        //                          .waitrequest
		.av_write                 (camera_dma_controller_avalon_dma_master_write),                                              //                          .write
		.av_writedata             (camera_dma_controller_avalon_dma_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                                       //               (terminated)
		.av_byteenable            (2'b11),                                                                                      //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                       //               (terminated)
		.av_begintransfer         (1'b0),                                                                                       //               (terminated)
		.av_chipselect            (1'b0),                                                                                       //               (terminated)
		.av_read                  (1'b0),                                                                                       //               (terminated)
		.av_readdata              (),                                                                                           //               (terminated)
		.av_readdatavalid         (),                                                                                           //               (terminated)
		.av_lock                  (1'b0),                                                                                       //               (terminated)
		.av_debugaccess           (1'b0),                                                                                       //               (terminated)
		.uav_clken                (),                                                                                           //               (terminated)
		.av_clken                 (1'b1),                                                                                       //               (terminated)
		.uav_response             (2'b00),                                                                                      //               (terminated)
		.av_response              (),                                                                                           //               (terminated)
		.uav_writeresponserequest (),                                                                                           //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                       //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                       //               (terminated)
		.av_writeresponsevalid    ()                                                                                            //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) lcd_dma_controller_avalon_dma_master_translator (
		.clk                      (sys_clk),                                                                                 //                       clk.clk
		.reset                    (cpu_jtag_debug_module_reset_reset),                                                       //                     reset.reset
		.uav_address              (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (lcd_dma_controller_avalon_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (lcd_dma_controller_avalon_dma_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (lcd_dma_controller_avalon_dma_master_read),                                               //                          .read
		.av_readdata              (lcd_dma_controller_avalon_dma_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (lcd_dma_controller_avalon_dma_master_readdatavalid),                                      //                          .readdatavalid
		.av_lock                  (lcd_dma_controller_avalon_dma_master_lock),                                               //                          .lock
		.av_burstcount            (1'b1),                                                                                    //               (terminated)
		.av_byteenable            (2'b11),                                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                    //               (terminated)
		.av_begintransfer         (1'b0),                                                                                    //               (terminated)
		.av_chipselect            (1'b0),                                                                                    //               (terminated)
		.av_write                 (1'b0),                                                                                    //               (terminated)
		.av_writedata             (16'b0000000000000000),                                                                    //               (terminated)
		.av_debugaccess           (1'b0),                                                                                    //               (terminated)
		.uav_clken                (),                                                                                        //               (terminated)
		.av_clken                 (1'b1),                                                                                    //               (terminated)
		.uav_response             (2'b00),                                                                                   //               (terminated)
		.av_response              (),                                                                                        //               (terminated)
		.uav_writeresponserequest (),                                                                                        //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                    //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                    //               (terminated)
		.av_writeresponsevalid    ()                                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) vga_dma_controller_avalon_dma_master_translator (
		.clk                      (sys_clk),                                                                                 //                       clk.clk
		.reset                    (cpu_jtag_debug_module_reset_reset),                                                       //                     reset.reset
		.uav_address              (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (vga_dma_controller_avalon_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (vga_dma_controller_avalon_dma_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (vga_dma_controller_avalon_dma_master_read),                                               //                          .read
		.av_readdata              (vga_dma_controller_avalon_dma_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (vga_dma_controller_avalon_dma_master_readdatavalid),                                      //                          .readdatavalid
		.av_lock                  (vga_dma_controller_avalon_dma_master_lock),                                               //                          .lock
		.av_burstcount            (1'b1),                                                                                    //               (terminated)
		.av_byteenable            (2'b11),                                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                    //               (terminated)
		.av_begintransfer         (1'b0),                                                                                    //               (terminated)
		.av_chipselect            (1'b0),                                                                                    //               (terminated)
		.av_write                 (1'b0),                                                                                    //               (terminated)
		.av_writedata             (16'b0000000000000000),                                                                    //               (terminated)
		.av_debugaccess           (1'b0),                                                                                    //               (terminated)
		.uav_clken                (),                                                                                        //               (terminated)
		.av_clken                 (1'b1),                                                                                    //               (terminated)
		.uav_response             (2'b00),                                                                                   //               (terminated)
		.av_response              (),                                                                                        //               (terminated)
		.uav_writeresponserequest (),                                                                                        //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                    //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                    //               (terminated)
		.av_writeresponsevalid    ()                                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) videoconferencing_dma_0_avalon_master_translator (
		.clk                      (sys_clk),                                                                                  //                       clk.clk
		.reset                    (rst_controller_006_reset_out_reset),                                                       //                     reset.reset
		.uav_address              (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (videoconferencing_dma_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (videoconferencing_dma_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (videoconferencing_dma_0_avalon_master_byteenable),                                         //                          .byteenable
		.av_write                 (videoconferencing_dma_0_avalon_master_write),                                              //                          .write
		.av_writedata             (videoconferencing_dma_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                                     //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                     //               (terminated)
		.av_begintransfer         (1'b0),                                                                                     //               (terminated)
		.av_chipselect            (1'b0),                                                                                     //               (terminated)
		.av_read                  (1'b0),                                                                                     //               (terminated)
		.av_readdata              (),                                                                                         //               (terminated)
		.av_readdatavalid         (),                                                                                         //               (terminated)
		.av_lock                  (1'b0),                                                                                     //               (terminated)
		.av_debugaccess           (1'b0),                                                                                     //               (terminated)
		.uav_clken                (),                                                                                         //               (terminated)
		.av_clken                 (1'b1),                                                                                     //               (terminated)
		.uav_response             (2'b00),                                                                                    //               (terminated)
		.av_response              (),                                                                                         //               (terminated)
		.uav_writeresponserequest (),                                                                                         //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                     //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                     //               (terminated)
		.av_writeresponsevalid    ()                                                                                          //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                      (sys_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_chipselect            (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (sys_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (21),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) flash_flash_data_translator (
		.clk                      (sys_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                          //                    reset.reset
		.uav_address              (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (flash_flash_data_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (flash_flash_data_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (flash_flash_data_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (flash_flash_data_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (flash_flash_data_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (flash_flash_data_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (flash_flash_data_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (flash_flash_data_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (sys_clk),                                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) interval_timer_s1_translator (
		.clk                      (sys_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address              (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (interval_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (interval_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (interval_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (interval_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (interval_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (sys_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) red_leds_avalon_parallel_port_slave_translator (
		.clk                      (sys_clk),                                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                 //                    reset.reset
		.uav_address              (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (red_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                                               //              (terminated)
		.av_burstcount            (),                                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                                               //              (terminated)
		.av_lock                  (),                                                                                               //              (terminated)
		.av_clken                 (),                                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                                           //              (terminated)
		.av_debugaccess           (),                                                                                               //              (terminated)
		.av_outputenable          (),                                                                                               //              (terminated)
		.uav_response             (),                                                                                               //              (terminated)
		.av_response              (2'b00),                                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) green_leds_avalon_parallel_port_slave_translator (
		.clk                      (sys_clk),                                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                   //                    reset.reset
		.uav_address              (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (green_leds_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                                 //              (terminated)
		.av_lock                  (),                                                                                                 //              (terminated)
		.av_clken                 (),                                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                                 //              (terminated)
		.uav_response             (),                                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex3_hex0_avalon_parallel_port_slave_translator (
		.clk                      (sys_clk),                                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                  //                    reset.reset
		.uav_address              (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (hex3_hex0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                                //              (terminated)
		.av_burstcount            (),                                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                                //              (terminated)
		.av_lock                  (),                                                                                                //              (terminated)
		.av_clken                 (),                                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                                //              (terminated)
		.av_outputenable          (),                                                                                                //              (terminated)
		.uav_response             (),                                                                                                //              (terminated)
		.av_response              (2'b00),                                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex7_hex4_avalon_parallel_port_slave_translator (
		.clk                      (sys_clk),                                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                  //                    reset.reset
		.uav_address              (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (hex7_hex4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                                //              (terminated)
		.av_burstcount            (),                                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                                //              (terminated)
		.av_lock                  (),                                                                                                //              (terminated)
		.av_clken                 (),                                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                                //              (terminated)
		.av_outputenable          (),                                                                                                //              (terminated)
		.uav_response             (),                                                                                                //              (terminated)
		.av_response              (2'b00),                                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) slider_switches_avalon_parallel_port_slave_translator (
		.clk                      (sys_clk),                                                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                        //                    reset.reset
		.uav_address              (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (slider_switches_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                                      //              (terminated)
		.av_lock                  (),                                                                                                      //              (terminated)
		.av_clken                 (),                                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                                      //              (terminated)
		.uav_response             (),                                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pushbuttons_avalon_parallel_port_slave_translator (
		.clk                      (sys_clk),                                                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                    //                    reset.reset
		.uav_address              (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (pushbuttons_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                                  //              (terminated)
		.av_lock                  (),                                                                                                  //              (terminated)
		.av_clken                 (),                                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                                  //              (terminated)
		.uav_response             (),                                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) expansion_jp5_avalon_parallel_port_slave_translator (
		.clk                      (sys_clk),                                                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                      //                    reset.reset
		.uav_address              (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (expansion_jp5_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                                    //              (terminated)
		.av_lock                  (),                                                                                                    //              (terminated)
		.av_clken                 (),                                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                                    //              (terminated)
		.uav_response             (),                                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) serial_port_avalon_rs232_slave_translator (
		.clk                      (sys_clk),                                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (serial_port_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_debugaccess           (),                                                                                          //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) char_lcd_16x2_avalon_lcd_slave_translator (
		.clk                      (sys_clk),                                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (char_lcd_16x2_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_byteenable            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_debugaccess           (),                                                                                          //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ps2_port_avalon_ps2_slave_translator (
		.clk                      (sys_clk),                                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (ps2_port_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                                     //              (terminated)
		.av_lock                  (),                                                                                     //              (terminated)
		.av_clken                 (),                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                 //              (terminated)
		.av_debugaccess           (),                                                                                     //              (terminated)
		.av_outputenable          (),                                                                                     //              (terminated)
		.uav_response             (),                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (20),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sram_avalon_sram_slave_translator (
		.clk                      (sys_clk),                                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sram_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sram_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sram_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sram_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sram_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sram_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_chipselect            (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) vga_char_buffer_avalon_char_control_slave_translator (
		.clk                      (sys_clk),                                                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                       //                    reset.reset
		.uav_address              (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (vga_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                                                     //              (terminated)
		.av_lock                  (),                                                                                                     //              (terminated)
		.av_clken                 (),                                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                                 //              (terminated)
		.av_debugaccess           (),                                                                                                     //              (terminated)
		.av_outputenable          (),                                                                                                     //              (terminated)
		.uav_response             (),                                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) vga_char_buffer_avalon_char_buffer_slave_translator (
		.clk                      (sys_clk),                                                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                      //                    reset.reset
		.uav_address              (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                                    //              (terminated)
		.av_lock                  (),                                                                                                    //              (terminated)
		.av_clken                 (),                                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                                    //              (terminated)
		.uav_response             (),                                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onboard_av_avalon_av_config_slave_translator (
		.clk                      (sys_clk),                                                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                               //                    reset.reset
		.uav_address              (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (onboard_av_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer         (),                                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                                             //              (terminated)
		.av_burstcount            (),                                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                                             //              (terminated)
		.av_lock                  (),                                                                                             //              (terminated)
		.av_chipselect            (),                                                                                             //              (terminated)
		.av_clken                 (),                                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                                         //              (terminated)
		.av_debugaccess           (),                                                                                             //              (terminated)
		.av_outputenable          (),                                                                                             //              (terminated)
		.uav_response             (),                                                                                             //              (terminated)
		.av_response              (2'b00),                                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ps2_port_dual_avalon_ps2_slave_translator (
		.clk                      (sys_clk),                                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (ps2_port_dual_avalon_ps2_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_debugaccess           (),                                                                                          //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_avalon_audio_slave_translator (
		.clk                      (sys_clk),                                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address              (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_avalon_audio_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_avalon_audio_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (audio_avalon_audio_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (audio_avalon_audio_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_avalon_audio_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (audio_avalon_audio_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_byteenable            (),                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) flash_flash_erase_control_translator (
		.clk                      (sys_clk),                                                                              //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (flash_flash_erase_control_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read                  (flash_flash_erase_control_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (flash_flash_erase_control_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (flash_flash_erase_control_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (flash_flash_erase_control_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (flash_flash_erase_control_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (flash_flash_erase_control_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_address               (),                                                                                     //              (terminated)
		.av_begintransfer         (),                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                                     //              (terminated)
		.av_lock                  (),                                                                                     //              (terminated)
		.av_clken                 (),                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                 //              (terminated)
		.av_debugaccess           (),                                                                                     //              (terminated)
		.av_outputenable          (),                                                                                     //              (terminated)
		.uav_response             (),                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_card_avalon_sdcard_slave_translator (
		.clk                      (sys_clk),                                                                                //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sd_card_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) irda_avalon_irda_slave_translator (
		.clk                      (sys_clk),                                                                           //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                                //                    reset.reset
		.uav_address              (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (irda_avalon_irda_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (irda_avalon_irda_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (irda_avalon_irda_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (irda_avalon_irda_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (irda_avalon_irda_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (irda_avalon_irda_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (irda_avalon_irda_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) video_in_dma_controller_avalon_dma_control_slave_translator (
		.clk                      (sys_clk),                                                                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                              //                    reset.reset
		.uav_address              (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer         (),                                                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                                                            //              (terminated)
		.av_burstcount            (),                                                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                                                            //              (terminated)
		.av_lock                  (),                                                                                                            //              (terminated)
		.av_chipselect            (),                                                                                                            //              (terminated)
		.av_clken                 (),                                                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                                                        //              (terminated)
		.av_debugaccess           (),                                                                                                            //              (terminated)
		.av_outputenable          (),                                                                                                            //              (terminated)
		.uav_response             (),                                                                                                            //              (terminated)
		.av_response              (2'b00),                                                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) camera_dma_controller_avalon_dma_control_slave_translator (
		.clk                      (sys_clk),                                                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                            //                    reset.reset
		.uav_address              (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (camera_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer         (),                                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                                          //              (terminated)
		.av_lock                  (),                                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                                          //              (terminated)
		.av_clken                 (),                                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                                      //              (terminated)
		.av_debugaccess           (),                                                                                                          //              (terminated)
		.av_outputenable          (),                                                                                                          //              (terminated)
		.uav_response             (),                                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) camera_config_avalon_av_config_slave_translator (
		.clk                      (sys_clk),                                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                  //                    reset.reset
		.uav_address              (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (camera_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer         (),                                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                                //              (terminated)
		.av_burstcount            (),                                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                                //              (terminated)
		.av_lock                  (),                                                                                                //              (terminated)
		.av_chipselect            (),                                                                                                //              (terminated)
		.av_clken                 (),                                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                                //              (terminated)
		.av_outputenable          (),                                                                                                //              (terminated)
		.uav_response             (),                                                                                                //              (terminated)
		.av_response              (2'b00),                                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) accelerometer_avalon_accelerometer_spi_mode_slave_translator (
		.clk                      (sys_clk),                                                                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                               //                    reset.reset
		.uav_address              (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer         (),                                                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                                                             //              (terminated)
		.av_burstcount            (),                                                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                                                             //              (terminated)
		.av_lock                  (),                                                                                                             //              (terminated)
		.av_chipselect            (),                                                                                                             //              (terminated)
		.av_clken                 (),                                                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                                                         //              (terminated)
		.av_debugaccess           (),                                                                                                             //              (terminated)
		.av_outputenable          (),                                                                                                             //              (terminated)
		.uav_response             (),                                                                                                             //              (terminated)
		.av_response              (2'b00),                                                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (5),
		.AV_WRITE_WAIT_CYCLES           (5),
		.AV_SETUP_WAIT_CYCLES           (5),
		.AV_DATA_HOLD_CYCLES            (5)
	) usb_avalon_usb_slave_translator (
		.clk                      (sys_clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address              (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (usb_avalon_usb_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (usb_avalon_usb_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (usb_avalon_usb_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (usb_avalon_usb_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (usb_avalon_usb_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (usb_avalon_usb_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                //              (terminated)
		.av_burstcount            (),                                                                                //              (terminated)
		.av_byteenable            (),                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                //              (terminated)
		.av_lock                  (),                                                                                //              (terminated)
		.av_clken                 (),                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                //              (terminated)
		.uav_response             (),                                                                                //              (terminated)
		.av_response              (2'b00),                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_char_buffer_avalon_char_control_slave_translator (
		.clk                      (sys_clk),                                                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                       //                    reset.reset
		.uav_address              (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (lcd_char_buffer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                                                     //              (terminated)
		.av_lock                  (),                                                                                                     //              (terminated)
		.av_clken                 (),                                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                                 //              (terminated)
		.av_debugaccess           (),                                                                                                     //              (terminated)
		.av_outputenable          (),                                                                                                     //              (terminated)
		.uav_response             (),                                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_char_buffer_avalon_char_buffer_slave_translator (
		.clk                      (sys_clk),                                                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                      //                    reset.reset
		.uav_address              (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                                    //              (terminated)
		.av_lock                  (),                                                                                                    //              (terminated)
		.av_clken                 (),                                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                                    //              (terminated)
		.uav_response             (),                                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) enet_control_port_translator (
		.clk                      (sys_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_005_reset_out_reset),                                           //                    reset.reset
		.uav_address              (enet_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (enet_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (enet_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (enet_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (enet_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (enet_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (enet_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (enet_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (enet_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (enet_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (enet_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (enet_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (enet_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (enet_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (enet_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (enet_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (enet_control_port_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_chipselect            (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) packet_memory_s1_translator (
		.clk                      (sys_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_005_reset_out_reset),                                          //                    reset.reset
		.uav_address              (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (packet_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (packet_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (packet_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (packet_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (packet_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (packet_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (packet_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) descriptor_memory_s1_translator (
		.clk                      (sys_clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_005_reset_out_reset),                                              //                    reset.reset
		.uav_address              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (descriptor_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (descriptor_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                                //              (terminated)
		.av_begintransfer         (),                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                //              (terminated)
		.av_burstcount            (),                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                //              (terminated)
		.av_lock                  (),                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                //              (terminated)
		.uav_response             (),                                                                                //              (terminated)
		.av_response              (2'b00),                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_dma_controller_avalon_dma_control_slave_translator (
		.clk                      (sys_clk),                                                                                                //                      clk.clk
		.reset                    (cpu_jtag_debug_module_reset_reset),                                                                      //                    reset.reset
		.uav_address              (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer         (),                                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                                       //              (terminated)
		.av_lock                  (),                                                                                                       //              (terminated)
		.av_chipselect            (),                                                                                                       //              (terminated)
		.av_clken                 (),                                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                                       //              (terminated)
		.uav_response             (),                                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) vga_dma_controller_avalon_dma_control_slave_translator (
		.clk                      (sys_clk),                                                                                                //                      clk.clk
		.reset                    (cpu_jtag_debug_module_reset_reset),                                                                      //                    reset.reset
		.uav_address              (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (vga_dma_controller_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer         (),                                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                                       //              (terminated)
		.av_lock                  (),                                                                                                       //              (terminated)
		.av_chipselect            (),                                                                                                       //              (terminated)
		.av_clken                 (),                                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                                       //              (terminated)
		.uav_response             (),                                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) videoconferencing_dma_0_avalon_slave_translator (
		.clk                      (sys_clk),                                                                                         //                      clk.clk
		.reset                    (rst_controller_006_reset_out_reset),                                                              //                    reset.reset
		.uav_address              (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (videoconferencing_dma_0_avalon_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                                //              (terminated)
		.av_burstcount            (),                                                                                                //              (terminated)
		.av_byteenable            (),                                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                                //              (terminated)
		.av_lock                  (),                                                                                                //              (terminated)
		.av_clken                 (),                                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                                //              (terminated)
		.av_outputenable          (),                                                                                                //              (terminated)
		.uav_response             (),                                                                                                //              (terminated)
		.av_response              (2'b00),                                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                             //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_THREAD_ID_H           (101),
		.PKT_THREAD_ID_L           (101),
		.PKT_CACHE_H               (108),
		.PKT_CACHE_L               (105),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.ST_DATA_W                 (111),
		.ST_CHANNEL_W              (38),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (sys_clk),                                                                            //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                               //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                              //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_THREAD_ID_H           (101),
		.PKT_THREAD_ID_L           (101),
		.PKT_CACHE_H               (108),
		.PKT_CACHE_L               (105),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.ST_DATA_W                 (111),
		.ST_CHANNEL_W              (38),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (sys_clk),                                                                     //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address              (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                  //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                   //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                          //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                            //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                  //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (77),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (38),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (6),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent (
		.clk                     (sys_clk),                                                                                               //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.av_address              (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_016_src1_valid),                                                                         //        rp.valid
		.rp_data                 (rsp_xbar_demux_016_src1_data),                                                                          //          .data
		.rp_channel              (rsp_xbar_demux_016_src1_channel),                                                                       //          .channel
		.rp_startofpacket        (rsp_xbar_demux_016_src1_startofpacket),                                                                 //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_016_src1_endofpacket),                                                                   //          .endofpacket
		.rp_ready                (rsp_xbar_demux_016_src1_ready),                                                                         //          .ready
		.av_response             (),                                                                                                      // (terminated)
		.av_writeresponserequest (1'b0),                                                                                                  // (terminated)
		.av_writeresponsevalid   ()                                                                                                       // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (77),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (38),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent (
		.clk                     (sys_clk),                                                                                             //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.av_address              (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_016_src2_valid),                                                                       //        rp.valid
		.rp_data                 (rsp_xbar_demux_016_src2_data),                                                                        //          .data
		.rp_channel              (rsp_xbar_demux_016_src2_channel),                                                                     //          .channel
		.rp_startofpacket        (rsp_xbar_demux_016_src2_startofpacket),                                                               //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_016_src2_endofpacket),                                                                 //          .endofpacket
		.rp_ready                (rsp_xbar_demux_016_src2_ready),                                                                       //          .ready
		.av_response             (),                                                                                                    // (terminated)
		.av_writeresponserequest (1'b0),                                                                                                // (terminated)
		.av_writeresponsevalid   ()                                                                                                     // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (77),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (38),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent (
		.clk                     (sys_clk),                                                                                          //       clk.clk
		.reset                   (cpu_jtag_debug_module_reset_reset),                                                                // clk_reset.reset
		.av_address              (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_016_src3_valid),                                                                    //        rp.valid
		.rp_data                 (rsp_xbar_demux_016_src3_data),                                                                     //          .data
		.rp_channel              (rsp_xbar_demux_016_src3_channel),                                                                  //          .channel
		.rp_startofpacket        (rsp_xbar_demux_016_src3_startofpacket),                                                            //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_016_src3_endofpacket),                                                              //          .endofpacket
		.rp_ready                (rsp_xbar_demux_016_src3_ready),                                                                    //          .ready
		.av_response             (),                                                                                                 // (terminated)
		.av_writeresponserequest (1'b0),                                                                                             // (terminated)
		.av_writeresponsevalid   ()                                                                                                  // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (77),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (38),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent (
		.clk                     (sys_clk),                                                                                          //       clk.clk
		.reset                   (cpu_jtag_debug_module_reset_reset),                                                                // clk_reset.reset
		.av_address              (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_016_src4_valid),                                                                    //        rp.valid
		.rp_data                 (rsp_xbar_demux_016_src4_data),                                                                     //          .data
		.rp_channel              (rsp_xbar_demux_016_src4_channel),                                                                  //          .channel
		.rp_startofpacket        (rsp_xbar_demux_016_src4_startofpacket),                                                            //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_016_src4_endofpacket),                                                              //          .endofpacket
		.rp_ready                (rsp_xbar_demux_016_src4_ready),                                                                    //          .ready
		.av_response             (),                                                                                                 // (terminated)
		.av_writeresponserequest (1'b0),                                                                                             // (terminated)
		.av_writeresponsevalid   ()                                                                                                  // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (77),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (38),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (5),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent (
		.clk                     (sys_clk),                                                                                           //       clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                                // clk_reset.reset
		.av_address              (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_016_src5_valid),                                                                     //        rp.valid
		.rp_data                 (rsp_xbar_demux_016_src5_data),                                                                      //          .data
		.rp_channel              (rsp_xbar_demux_016_src5_channel),                                                                   //          .channel
		.rp_startofpacket        (rsp_xbar_demux_016_src5_startofpacket),                                                             //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_016_src5_endofpacket),                                                               //          .endofpacket
		.rp_ready                (rsp_xbar_demux_016_src5_ready),                                                                     //          .ready
		.av_response             (),                                                                                                  // (terminated)
		.av_writeresponserequest (1'b0),                                                                                              // (terminated)
		.av_writeresponsevalid   ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                  //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) flash_flash_data_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (flash_flash_data_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (flash_flash_data_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (flash_flash_data_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (flash_flash_data_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (flash_flash_data_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (flash_flash_data_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                          //                .channel
		.rf_sink_ready           (flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (flash_flash_data_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (flash_flash_data_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (flash_flash_data_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (flash_flash_data_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (flash_flash_data_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (flash_flash_data_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                               //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (flash_flash_data_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (flash_flash_data_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) interval_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                        //                .channel
		.rf_sink_ready           (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                           //       clk_reset.reset
		.m0_address              (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                                          //                .channel
		.rf_sink_ready           (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                           // clk_reset.reset
		.in_data           (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                                     // (terminated)
		.csr_readdata      (),                                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                     // (terminated)
		.almost_full_data  (),                                                                                                         // (terminated)
		.almost_empty_data (),                                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                                     // (terminated)
		.out_empty         (),                                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                                     // (terminated)
		.out_error         (),                                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                                     // (terminated)
		.out_channel       ()                                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                                            //                .channel
		.rf_sink_ready           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                            //       clk_reset.reset
		.m0_address              (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                                           //                .channel
		.rf_sink_ready           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                            // clk_reset.reset
		.in_data           (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                            //       clk_reset.reset
		.m0_address              (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                                           //                .channel
		.rf_sink_ready           (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                            // clk_reset.reset
		.in_data           (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                  //       clk_reset.reset
		.m0_address              (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                                                //                .channel
		.rf_sink_ready           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                  // clk_reset.reset
		.in_data           (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                            // (terminated)
		.almost_full_data  (),                                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                                            // (terminated)
		.out_empty         (),                                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                                            // (terminated)
		.out_error         (),                                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                                            // (terminated)
		.out_channel       ()                                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                              //       clk_reset.reset
		.m0_address              (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                                            //                .channel
		.rf_sink_ready           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                              // clk_reset.reset
		.in_data           (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                                        // (terminated)
		.csr_readdata      (),                                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                        // (terminated)
		.almost_full_data  (),                                                                                                            // (terminated)
		.almost_empty_data (),                                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                                        // (terminated)
		.out_empty         (),                                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                                        // (terminated)
		.out_error         (),                                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                                        // (terminated)
		.out_channel       ()                                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                //       clk_reset.reset
		.m0_address              (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                                              //                .channel
		.rf_sink_ready           (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                // clk_reset.reset
		.in_data           (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                                          // (terminated)
		.csr_readdata      (),                                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                          // (terminated)
		.almost_full_data  (),                                                                                                              // (terminated)
		.almost_empty_data (),                                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                                          // (terminated)
		.out_empty         (),                                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                                          // (terminated)
		.out_error         (),                                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                                          // (terminated)
		.out_channel       ()                                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                                    //                .channel
		.rf_sink_ready           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                         //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                         //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                          //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                                       //                .channel
		.rf_sink_ready           (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                                               //                .channel
		.rf_sink_ready           (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                             //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                             //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                              //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                       //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                           //                .channel
		.rf_sink_ready           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (sys_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                                  // (terminated)
		.out_startofpacket (),                                                                                      // (terminated)
		.out_endofpacket   (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                 //       clk_reset.reset
		.m0_address              (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                                                               //                .channel
		.rf_sink_ready           (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                 // clk_reset.reset
		.in_data           (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                                           // (terminated)
		.csr_readdata      (),                                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                           // (terminated)
		.almost_full_data  (),                                                                                                               // (terminated)
		.almost_empty_data (),                                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                                           // (terminated)
		.out_empty         (),                                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                                           // (terminated)
		.out_error         (),                                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                                           // (terminated)
		.out_channel       ()                                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                //       clk_reset.reset
		.m0_address              (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                                               //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                                               //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                                                //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                                         //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                                             //                .channel
		.rf_sink_ready           (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                // clk_reset.reset
		.in_data           (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                                          // (terminated)
		.csr_readdata      (),                                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                          // (terminated)
		.almost_full_data  (),                                                                                                              // (terminated)
		.almost_empty_data (),                                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                                          // (terminated)
		.out_empty         (),                                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                                          // (terminated)
		.out_error         (),                                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                                          // (terminated)
		.out_channel       ()                                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src19_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src19_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src19_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src19_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src19_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src19_channel),                                                                       //                .channel
		.rf_sink_ready           (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src20_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src20_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src20_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src20_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src20_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src20_channel),                                                                    //                .channel
		.rf_sink_ready           (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src21_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src21_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src21_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src21_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src21_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src21_channel),                                                              //                .channel
		.rf_sink_ready           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) flash_flash_erase_control_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src22_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src22_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src22_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src22_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src22_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src22_channel),                                                               //                .channel
		.rf_sink_ready           (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src23_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src23_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src23_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src23_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src23_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src23_channel),                                                                 //                .channel
		.rf_sink_ready           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src24_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src24_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src24_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src24_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src24_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src24_channel),                                                            //                .channel
		.rf_sink_ready           (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                        //       clk_reset.reset
		.m0_address              (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src25_ready),                                                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src25_valid),                                                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_001_src25_data),                                                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src25_startofpacket),                                                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src25_endofpacket),                                                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src25_channel),                                                                                      //                .channel
		.rf_sink_ready           (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                        // clk_reset.reset
		.in_data           (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                  // (terminated)
		.almost_full_data  (),                                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                                  // (terminated)
		.out_empty         (),                                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                                  // (terminated)
		.out_error         (),                                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                                  // (terminated)
		.out_channel       ()                                                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                      //       clk_reset.reset
		.m0_address              (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src26_ready),                                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src26_valid),                                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src26_data),                                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src26_startofpacket),                                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src26_endofpacket),                                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src26_channel),                                                                                    //                .channel
		.rf_sink_ready           (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                      // clk_reset.reset
		.in_data           (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                // (terminated)
		.almost_full_data  (),                                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                                // (terminated)
		.out_empty         (),                                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                                // (terminated)
		.out_error         (),                                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                                // (terminated)
		.out_channel       ()                                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                            //       clk_reset.reset
		.m0_address              (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src27_ready),                                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src27_valid),                                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src27_data),                                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src27_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src27_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src27_channel),                                                                          //                .channel
		.rf_sink_ready           (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                            // clk_reset.reset
		.in_data           (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                         //       clk_reset.reset
		.m0_address              (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                                                        //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                                                        //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                                                         //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                                                  //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                                                      //                .channel
		.rf_sink_ready           (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                         // clk_reset.reset
		.in_data           (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                   // (terminated)
		.almost_full_data  (),                                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                                   // (terminated)
		.out_empty         (),                                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                                   // (terminated)
		.out_error         (),                                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                                   // (terminated)
		.out_channel       ()                                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src29_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src29_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src29_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src29_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src29_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src29_channel),                                                          //                .channel
		.rf_sink_ready           (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                 //       clk_reset.reset
		.m0_address              (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src30_ready),                                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src30_valid),                                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src30_data),                                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src30_startofpacket),                                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src30_endofpacket),                                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src30_channel),                                                                               //                .channel
		.rf_sink_ready           (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                 // clk_reset.reset
		.in_data           (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                                           // (terminated)
		.csr_readdata      (),                                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                           // (terminated)
		.almost_full_data  (),                                                                                                               // (terminated)
		.almost_empty_data (),                                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                                           // (terminated)
		.out_empty         (),                                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                                           // (terminated)
		.out_error         (),                                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                                           // (terminated)
		.out_channel       ()                                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (67),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (73),
		.PKT_DEST_ID_L             (68),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (77),
		.PKT_PROTECTION_L          (75),
		.PKT_RESPONSE_STATUS_H     (83),
		.PKT_RESPONSE_STATUS_L     (82),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                //       clk_reset.reset
		.m0_address              (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_004_source0_ready),                                                                               //              cp.ready
		.cp_valid                (burst_adapter_004_source0_valid),                                                                               //                .valid
		.cp_data                 (burst_adapter_004_source0_data),                                                                                //                .data
		.cp_startofpacket        (burst_adapter_004_source0_startofpacket),                                                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_004_source0_endofpacket),                                                                         //                .endofpacket
		.cp_channel              (burst_adapter_004_source0_channel),                                                                             //                .channel
		.rf_sink_ready           (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                // clk_reset.reset
		.in_data           (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                                          // (terminated)
		.csr_readdata      (),                                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                          // (terminated)
		.almost_full_data  (),                                                                                                              // (terminated)
		.almost_empty_data (),                                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                                          // (terminated)
		.out_empty         (),                                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                                          // (terminated)
		.out_error         (),                                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                                          // (terminated)
		.out_channel       ()                                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) enet_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (enet_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (enet_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (enet_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (enet_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (enet_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (enet_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (enet_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (enet_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (enet_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (enet_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (enet_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (enet_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (enet_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (enet_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (enet_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (enet_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src32_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src32_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src32_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src32_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src32_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src32_channel),                                                       //                .channel
		.rf_sink_ready           (enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (enet_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (enet_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (enet_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (enet_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (enet_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (enet_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (enet_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (enet_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) packet_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (packet_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src33_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src33_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_001_src33_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src33_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src33_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src33_channel),                                                      //                .channel
		.rf_sink_ready           (packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (packet_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (packet_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (packet_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (packet_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (packet_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (packet_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                               //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (packet_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (packet_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src34_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src34_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src34_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src34_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src34_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src34_channel),                                                          //                .channel
		.rf_sink_ready           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_005_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                          //             clk.clk
		.reset                   (cpu_jtag_debug_module_reset_reset),                                                                                //       clk_reset.reset
		.m0_address              (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src35_ready),                                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src35_valid),                                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src35_data),                                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src35_startofpacket),                                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src35_endofpacket),                                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src35_channel),                                                                                 //                .channel
		.rf_sink_ready           (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                          //       clk.clk
		.reset             (cpu_jtag_debug_module_reset_reset),                                                                                // clk_reset.reset
		.in_data           (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                             // (terminated)
		.almost_full_data  (),                                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                                             // (terminated)
		.out_empty         (),                                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                                             // (terminated)
		.out_error         (),                                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                                             // (terminated)
		.out_channel       ()                                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                          //             clk.clk
		.reset                   (cpu_jtag_debug_module_reset_reset),                                                                                //       clk_reset.reset
		.m0_address              (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src36_ready),                                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src36_valid),                                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src36_data),                                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src36_startofpacket),                                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src36_endofpacket),                                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src36_channel),                                                                                 //                .channel
		.rf_sink_ready           (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                          //       clk.clk
		.reset             (cpu_jtag_debug_module_reset_reset),                                                                                // clk_reset.reset
		.in_data           (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                             // (terminated)
		.almost_full_data  (),                                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                                             // (terminated)
		.out_empty         (),                                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                                             // (terminated)
		.out_error         (),                                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                                             // (terminated)
		.out_channel       ()                                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (104),
		.PKT_PROTECTION_L          (102),
		.PKT_RESPONSE_STATUS_H     (110),
		.PKT_RESPONSE_STATUS_L     (109),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (38),
		.ST_DATA_W                 (111),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (sys_clk),                                                                                                   //             clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src37_ready),                                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src37_valid),                                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src37_data),                                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src37_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src37_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src37_channel),                                                                          //                .channel
		.rf_sink_ready           (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (112),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sys_clk),                                                                                                   //       clk.clk
		.reset             (rst_controller_006_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	nios_system_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	nios_system_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                              //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_002 (
		.sink_ready         (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (video_in_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                                             //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                                             //          .valid
		.src_data           (addr_router_002_src_data),                                                                              //          .data
		.src_channel        (addr_router_002_src_channel),                                                                           //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                                     //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                                        //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_003 (
		.sink_ready         (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (camera_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                                           //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                                           //          .valid
		.src_data           (addr_router_003_src_data),                                                                            //          .data
		.src_channel        (addr_router_003_src_channel),                                                                         //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                                   //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                                      //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_004 (
		.sink_ready         (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                          //       clk.clk
		.reset              (cpu_jtag_debug_module_reset_reset),                                                                // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                                        //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                                        //          .valid
		.src_data           (addr_router_004_src_data),                                                                         //          .data
		.src_channel        (addr_router_004_src_channel),                                                                      //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                                   //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_005 (
		.sink_ready         (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (vga_dma_controller_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                          //       clk.clk
		.reset              (cpu_jtag_debug_module_reset_reset),                                                                // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                                        //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                                        //          .valid
		.src_data           (addr_router_005_src_data),                                                                         //          .data
		.src_channel        (addr_router_005_src_channel),                                                                      //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                                   //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_006 (
		.sink_ready         (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (videoconferencing_dma_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                           //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                                                // clk_reset.reset
		.src_ready          (addr_router_006_src_ready),                                                                         //       src.ready
		.src_valid          (addr_router_006_src_valid),                                                                         //          .valid
		.src_data           (addr_router_006_src_data),                                                                          //          .data
		.src_channel        (addr_router_006_src_channel),                                                                       //          .channel
		.src_startofpacket  (addr_router_006_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (addr_router_006_src_endofpacket)                                                                    //          .endofpacket
	);

	nios_system_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	nios_system_id_router id_router_001 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                             //       src.ready
		.src_valid          (id_router_001_src_valid),                                             //          .valid
		.src_data           (id_router_001_src_data),                                              //          .data
		.src_channel        (id_router_001_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router id_router_002 (
		.sink_ready         (flash_flash_data_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (flash_flash_data_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (flash_flash_data_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (flash_flash_data_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (flash_flash_data_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                     //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                     //       src.ready
		.src_valid          (id_router_002_src_valid),                                                     //          .valid
		.src_data           (id_router_002_src_data),                                                      //          .data
		.src_channel        (id_router_002_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                //          .endofpacket
	);

	nios_system_id_router_003 id_router_003 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                //          .valid
		.src_data           (id_router_003_src_data),                                                                 //          .data
		.src_channel        (id_router_003_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                           //          .endofpacket
	);

	nios_system_id_router_003 id_router_004 (
		.sink_ready         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                      //       src.ready
		.src_valid          (id_router_004_src_valid),                                                      //          .valid
		.src_data           (id_router_004_src_data),                                                       //          .data
		.src_channel        (id_router_004_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                 //          .endofpacket
	);

	nios_system_id_router_003 id_router_005 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                        //       src.ready
		.src_valid          (id_router_005_src_valid),                                                        //          .valid
		.src_data           (id_router_005_src_data),                                                         //          .data
		.src_channel        (id_router_005_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                   //          .endofpacket
	);

	nios_system_id_router_003 id_router_006 (
		.sink_ready         (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (red_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                        //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                        //          .valid
		.src_data           (id_router_006_src_data),                                                                         //          .data
		.src_channel        (id_router_006_src_channel),                                                                      //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                                   //          .endofpacket
	);

	nios_system_id_router_003 id_router_007 (
		.sink_ready         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (green_leds_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                          //          .valid
		.src_data           (id_router_007_src_data),                                                                           //          .data
		.src_channel        (id_router_007_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_id_router_003 id_router_008 (
		.sink_ready         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex3_hex0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                         //          .valid
		.src_data           (id_router_008_src_data),                                                                          //          .data
		.src_channel        (id_router_008_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                    //          .endofpacket
	);

	nios_system_id_router_003 id_router_009 (
		.sink_ready         (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex7_hex4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_009_src_valid),                                                                         //          .valid
		.src_data           (id_router_009_src_data),                                                                          //          .data
		.src_channel        (id_router_009_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                                    //          .endofpacket
	);

	nios_system_id_router_003 id_router_010 (
		.sink_ready         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slider_switches_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                                                               //          .valid
		.src_data           (id_router_010_src_data),                                                                                //          .data
		.src_channel        (id_router_010_src_channel),                                                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                                          //          .endofpacket
	);

	nios_system_id_router_003 id_router_011 (
		.sink_ready         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pushbuttons_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                                           //       src.ready
		.src_valid          (id_router_011_src_valid),                                                                           //          .valid
		.src_data           (id_router_011_src_data),                                                                            //          .data
		.src_channel        (id_router_011_src_channel),                                                                         //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                                   //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                                      //          .endofpacket
	);

	nios_system_id_router_003 id_router_012 (
		.sink_ready         (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (expansion_jp5_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                                             //       src.ready
		.src_valid          (id_router_012_src_valid),                                                                             //          .valid
		.src_data           (id_router_012_src_data),                                                                              //          .data
		.src_channel        (id_router_012_src_channel),                                                                           //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                                                     //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                                        //          .endofpacket
	);

	nios_system_id_router_003 id_router_013 (
		.sink_ready         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (serial_port_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_013_src_valid),                                                                   //          .valid
		.src_data           (id_router_013_src_data),                                                                    //          .data
		.src_channel        (id_router_013_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                              //          .endofpacket
	);

	nios_system_id_router_014 id_router_014 (
		.sink_ready         (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (char_lcd_16x2_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_014_src_valid),                                                                   //          .valid
		.src_data           (id_router_014_src_data),                                                                    //          .data
		.src_channel        (id_router_014_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                              //          .endofpacket
	);

	nios_system_id_router_003 id_router_015 (
		.sink_ready         (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ps2_port_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                              //       src.ready
		.src_valid          (id_router_015_src_valid),                                                              //          .valid
		.src_data           (id_router_015_src_data),                                                               //          .data
		.src_channel        (id_router_015_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                         //          .endofpacket
	);

	nios_system_id_router_016 id_router_016 (
		.sink_ready         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                           //       src.ready
		.src_valid          (id_router_016_src_valid),                                                           //          .valid
		.src_data           (id_router_016_src_data),                                                            //          .data
		.src_channel        (id_router_016_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                      //          .endofpacket
	);

	nios_system_id_router_003 id_router_017 (
		.sink_ready         (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (vga_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                                              //       src.ready
		.src_valid          (id_router_017_src_valid),                                                                              //          .valid
		.src_data           (id_router_017_src_data),                                                                               //          .data
		.src_channel        (id_router_017_src_channel),                                                                            //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                                         //          .endofpacket
	);

	nios_system_id_router_014 id_router_018 (
		.sink_ready         (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (vga_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                                             //       src.ready
		.src_valid          (id_router_018_src_valid),                                                                             //          .valid
		.src_data           (id_router_018_src_data),                                                                              //          .data
		.src_channel        (id_router_018_src_channel),                                                                           //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                                                     //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                                        //          .endofpacket
	);

	nios_system_id_router_003 id_router_019 (
		.sink_ready         (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onboard_av_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_019_src_valid),                                                                      //          .valid
		.src_data           (id_router_019_src_data),                                                                       //          .data
		.src_channel        (id_router_019_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                                                 //          .endofpacket
	);

	nios_system_id_router_003 id_router_020 (
		.sink_ready         (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ps2_port_dual_avalon_ps2_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_020_src_valid),                                                                   //          .valid
		.src_data           (id_router_020_src_data),                                                                    //          .data
		.src_channel        (id_router_020_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                                              //          .endofpacket
	);

	nios_system_id_router_003 id_router_021 (
		.sink_ready         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_avalon_audio_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                             //       src.ready
		.src_valid          (id_router_021_src_valid),                                                             //          .valid
		.src_data           (id_router_021_src_data),                                                              //          .data
		.src_channel        (id_router_021_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                                        //          .endofpacket
	);

	nios_system_id_router_003 id_router_022 (
		.sink_ready         (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (flash_flash_erase_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                              //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                                              //       src.ready
		.src_valid          (id_router_022_src_valid),                                                              //          .valid
		.src_data           (id_router_022_src_data),                                                               //          .data
		.src_channel        (id_router_022_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                                         //          .endofpacket
	);

	nios_system_id_router_003 id_router_023 (
		.sink_ready         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_card_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                                                //       src.ready
		.src_valid          (id_router_023_src_valid),                                                                //          .valid
		.src_data           (id_router_023_src_data),                                                                 //          .data
		.src_channel        (id_router_023_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                                           //          .endofpacket
	);

	nios_system_id_router_003 id_router_024 (
		.sink_ready         (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (irda_avalon_irda_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                           //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                                           //       src.ready
		.src_valid          (id_router_024_src_valid),                                                           //          .valid
		.src_data           (id_router_024_src_data),                                                            //          .data
		.src_channel        (id_router_024_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                                      //          .endofpacket
	);

	nios_system_id_router_003 id_router_025 (
		.sink_ready         (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (video_in_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                              // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                                                     //       src.ready
		.src_valid          (id_router_025_src_valid),                                                                                     //          .valid
		.src_data           (id_router_025_src_data),                                                                                      //          .data
		.src_channel        (id_router_025_src_channel),                                                                                   //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                                                             //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                                                                //          .endofpacket
	);

	nios_system_id_router_003 id_router_026 (
		.sink_ready         (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (camera_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                            // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                                                                   //       src.ready
		.src_valid          (id_router_026_src_valid),                                                                                   //          .valid
		.src_data           (id_router_026_src_data),                                                                                    //          .data
		.src_channel        (id_router_026_src_channel),                                                                                 //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                                                           //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                                                              //          .endofpacket
	);

	nios_system_id_router_003 id_router_027 (
		.sink_ready         (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (camera_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_027_src_valid),                                                                         //          .valid
		.src_data           (id_router_027_src_data),                                                                          //          .data
		.src_channel        (id_router_027_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                                                    //          .endofpacket
	);

	nios_system_id_router_014 id_router_028 (
		.sink_ready         (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (accelerometer_avalon_accelerometer_spi_mode_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                               // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                                                                      //       src.ready
		.src_valid          (id_router_028_src_valid),                                                                                      //          .valid
		.src_data           (id_router_028_src_data),                                                                                       //          .data
		.src_channel        (id_router_028_src_channel),                                                                                    //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                                                              //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                                                                 //          .endofpacket
	);

	nios_system_id_router_003 id_router_029 (
		.sink_ready         (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (usb_avalon_usb_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_029_src_ready),                                                         //       src.ready
		.src_valid          (id_router_029_src_valid),                                                         //          .valid
		.src_data           (id_router_029_src_data),                                                          //          .data
		.src_channel        (id_router_029_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_029_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_029_src_endofpacket)                                                    //          .endofpacket
	);

	nios_system_id_router_003 id_router_030 (
		.sink_ready         (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_char_buffer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.src_ready          (id_router_030_src_ready),                                                                              //       src.ready
		.src_valid          (id_router_030_src_valid),                                                                              //          .valid
		.src_data           (id_router_030_src_data),                                                                               //          .data
		.src_channel        (id_router_030_src_channel),                                                                            //          .channel
		.src_startofpacket  (id_router_030_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (id_router_030_src_endofpacket)                                                                         //          .endofpacket
	);

	nios_system_id_router_014 id_router_031 (
		.sink_ready         (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_char_buffer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.src_ready          (id_router_031_src_ready),                                                                             //       src.ready
		.src_valid          (id_router_031_src_valid),                                                                             //          .valid
		.src_data           (id_router_031_src_data),                                                                              //          .data
		.src_channel        (id_router_031_src_channel),                                                                           //          .channel
		.src_startofpacket  (id_router_031_src_startofpacket),                                                                     //          .startofpacket
		.src_endofpacket    (id_router_031_src_endofpacket)                                                                        //          .endofpacket
	);

	nios_system_id_router_003 id_router_032 (
		.sink_ready         (enet_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (enet_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (enet_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (enet_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (enet_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                      //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_032_src_ready),                                                      //       src.ready
		.src_valid          (id_router_032_src_valid),                                                      //          .valid
		.src_data           (id_router_032_src_data),                                                       //          .data
		.src_channel        (id_router_032_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_032_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_032_src_endofpacket)                                                 //          .endofpacket
	);

	nios_system_id_router_003 id_router_033 (
		.sink_ready         (packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (packet_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                     //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_033_src_ready),                                                     //       src.ready
		.src_valid          (id_router_033_src_valid),                                                     //          .valid
		.src_data           (id_router_033_src_data),                                                      //          .data
		.src_channel        (id_router_033_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_033_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_033_src_endofpacket)                                                //          .endofpacket
	);

	nios_system_id_router_003 id_router_034 (
		.sink_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                         //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_034_src_ready),                                                         //       src.ready
		.src_valid          (id_router_034_src_valid),                                                         //          .valid
		.src_data           (id_router_034_src_data),                                                          //          .data
		.src_channel        (id_router_034_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_034_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_034_src_endofpacket)                                                    //          .endofpacket
	);

	nios_system_id_router_003 id_router_035 (
		.sink_ready         (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                                //       clk.clk
		.reset              (cpu_jtag_debug_module_reset_reset),                                                                      // clk_reset.reset
		.src_ready          (id_router_035_src_ready),                                                                                //       src.ready
		.src_valid          (id_router_035_src_valid),                                                                                //          .valid
		.src_data           (id_router_035_src_data),                                                                                 //          .data
		.src_channel        (id_router_035_src_channel),                                                                              //          .channel
		.src_startofpacket  (id_router_035_src_startofpacket),                                                                        //          .startofpacket
		.src_endofpacket    (id_router_035_src_endofpacket)                                                                           //          .endofpacket
	);

	nios_system_id_router_003 id_router_036 (
		.sink_ready         (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (vga_dma_controller_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                                //       clk.clk
		.reset              (cpu_jtag_debug_module_reset_reset),                                                                      // clk_reset.reset
		.src_ready          (id_router_036_src_ready),                                                                                //       src.ready
		.src_valid          (id_router_036_src_valid),                                                                                //          .valid
		.src_data           (id_router_036_src_data),                                                                                 //          .data
		.src_channel        (id_router_036_src_channel),                                                                              //          .channel
		.src_startofpacket  (id_router_036_src_startofpacket),                                                                        //          .startofpacket
		.src_endofpacket    (id_router_036_src_endofpacket)                                                                           //          .endofpacket
	);

	nios_system_id_router_003 id_router_037 (
		.sink_ready         (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (videoconferencing_dma_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sys_clk),                                                                                         //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_037_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_037_src_valid),                                                                         //          .valid
		.src_data           (id_router_037_src_data),                                                                          //          .data
		.src_channel        (id_router_037_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_037_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_037_src_endofpacket)                                                                    //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (100),
		.PKT_DEST_ID_L             (95),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (111),
		.ST_CHANNEL_W              (38),
		.VALID_WIDTH               (38),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (sys_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (38),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter (
		.clk                   (sys_clk),                             //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (38),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_001 (
		.clk                   (sys_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_016_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_016_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_016_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_016_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_016_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_016_src_ready),              //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (38),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_002 (
		.clk                   (sys_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (38),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_003 (
		.clk                   (sys_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_003_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_003_src_data),              //          .data
		.sink0_channel         (width_adapter_003_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_003_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_003_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_003_src_ready),             //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (38),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_004 (
		.clk                   (sys_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_004_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_004_source0_data),          //          .data
		.source0_channel       (burst_adapter_004_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_004_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_004_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_004_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_n),                          // reset_in0.reset
		.reset_in1  (~reset_n),                          // reset_in1.reset
		.reset_in2  (cpu_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk        (sys_clk),                           //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req  (),                                  // (terminated)
		.reset_in3  (1'b0),                              // (terminated)
		.reset_in4  (1'b0),                              // (terminated)
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (~reset_n),                           // reset_in1.reset
		.reset_in2  (cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.clk        (vga_clk_out_clk_clk),                //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (4),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (~reset_n),                           // reset_in1.reset
		.reset_in2  (~reset_n),                           // reset_in2.reset
		.reset_in3  (cpu_jtag_debug_module_reset_reset),  // reset_in3.reset
		.clk        (clk),                                //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_003 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk        (sys_clk),                            //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_004 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.reset_in2  (~reset_n),                           // reset_in2.reset
		.clk        (external_clocks_vga_clk_33_clk),     //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller_005 (
		.reset_in0  (~reset_n),                               // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk        (sys_clk),                                //       clk.clk
		.reset_out  (rst_controller_005_reset_out_reset),     // reset_out.reset
		.reset_req  (rst_controller_005_reset_out_reset_req), //          .reset_req
		.reset_in2  (1'b0),                                   // (terminated)
		.reset_in3  (1'b0),                                   // (terminated)
		.reset_in4  (1'b0),                                   // (terminated)
		.reset_in5  (1'b0),                                   // (terminated)
		.reset_in6  (1'b0),                                   // (terminated)
		.reset_in7  (1'b0),                                   // (terminated)
		.reset_in8  (1'b0),                                   // (terminated)
		.reset_in9  (1'b0),                                   // (terminated)
		.reset_in10 (1'b0),                                   // (terminated)
		.reset_in11 (1'b0),                                   // (terminated)
		.reset_in12 (1'b0),                                   // (terminated)
		.reset_in13 (1'b0),                                   // (terminated)
		.reset_in14 (1'b0),                                   // (terminated)
		.reset_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_006 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.clk        (sys_clk),                            //       clk.clk
		.reset_out  (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (sys_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (sys_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_001_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_001_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_001_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_001_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_001_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_001_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_001_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_001_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_001_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_001_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_001_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_001_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_001_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_001_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_001_src22_endofpacket),   //          .endofpacket
		.src23_ready         (cmd_xbar_demux_001_src23_ready),         //     src23.ready
		.src23_valid         (cmd_xbar_demux_001_src23_valid),         //          .valid
		.src23_data          (cmd_xbar_demux_001_src23_data),          //          .data
		.src23_channel       (cmd_xbar_demux_001_src23_channel),       //          .channel
		.src23_startofpacket (cmd_xbar_demux_001_src23_startofpacket), //          .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_001_src23_endofpacket),   //          .endofpacket
		.src24_ready         (cmd_xbar_demux_001_src24_ready),         //     src24.ready
		.src24_valid         (cmd_xbar_demux_001_src24_valid),         //          .valid
		.src24_data          (cmd_xbar_demux_001_src24_data),          //          .data
		.src24_channel       (cmd_xbar_demux_001_src24_channel),       //          .channel
		.src24_startofpacket (cmd_xbar_demux_001_src24_startofpacket), //          .startofpacket
		.src24_endofpacket   (cmd_xbar_demux_001_src24_endofpacket),   //          .endofpacket
		.src25_ready         (cmd_xbar_demux_001_src25_ready),         //     src25.ready
		.src25_valid         (cmd_xbar_demux_001_src25_valid),         //          .valid
		.src25_data          (cmd_xbar_demux_001_src25_data),          //          .data
		.src25_channel       (cmd_xbar_demux_001_src25_channel),       //          .channel
		.src25_startofpacket (cmd_xbar_demux_001_src25_startofpacket), //          .startofpacket
		.src25_endofpacket   (cmd_xbar_demux_001_src25_endofpacket),   //          .endofpacket
		.src26_ready         (cmd_xbar_demux_001_src26_ready),         //     src26.ready
		.src26_valid         (cmd_xbar_demux_001_src26_valid),         //          .valid
		.src26_data          (cmd_xbar_demux_001_src26_data),          //          .data
		.src26_channel       (cmd_xbar_demux_001_src26_channel),       //          .channel
		.src26_startofpacket (cmd_xbar_demux_001_src26_startofpacket), //          .startofpacket
		.src26_endofpacket   (cmd_xbar_demux_001_src26_endofpacket),   //          .endofpacket
		.src27_ready         (cmd_xbar_demux_001_src27_ready),         //     src27.ready
		.src27_valid         (cmd_xbar_demux_001_src27_valid),         //          .valid
		.src27_data          (cmd_xbar_demux_001_src27_data),          //          .data
		.src27_channel       (cmd_xbar_demux_001_src27_channel),       //          .channel
		.src27_startofpacket (cmd_xbar_demux_001_src27_startofpacket), //          .startofpacket
		.src27_endofpacket   (cmd_xbar_demux_001_src27_endofpacket),   //          .endofpacket
		.src28_ready         (cmd_xbar_demux_001_src28_ready),         //     src28.ready
		.src28_valid         (cmd_xbar_demux_001_src28_valid),         //          .valid
		.src28_data          (cmd_xbar_demux_001_src28_data),          //          .data
		.src28_channel       (cmd_xbar_demux_001_src28_channel),       //          .channel
		.src28_startofpacket (cmd_xbar_demux_001_src28_startofpacket), //          .startofpacket
		.src28_endofpacket   (cmd_xbar_demux_001_src28_endofpacket),   //          .endofpacket
		.src29_ready         (cmd_xbar_demux_001_src29_ready),         //     src29.ready
		.src29_valid         (cmd_xbar_demux_001_src29_valid),         //          .valid
		.src29_data          (cmd_xbar_demux_001_src29_data),          //          .data
		.src29_channel       (cmd_xbar_demux_001_src29_channel),       //          .channel
		.src29_startofpacket (cmd_xbar_demux_001_src29_startofpacket), //          .startofpacket
		.src29_endofpacket   (cmd_xbar_demux_001_src29_endofpacket),   //          .endofpacket
		.src30_ready         (cmd_xbar_demux_001_src30_ready),         //     src30.ready
		.src30_valid         (cmd_xbar_demux_001_src30_valid),         //          .valid
		.src30_data          (cmd_xbar_demux_001_src30_data),          //          .data
		.src30_channel       (cmd_xbar_demux_001_src30_channel),       //          .channel
		.src30_startofpacket (cmd_xbar_demux_001_src30_startofpacket), //          .startofpacket
		.src30_endofpacket   (cmd_xbar_demux_001_src30_endofpacket),   //          .endofpacket
		.src31_ready         (cmd_xbar_demux_001_src31_ready),         //     src31.ready
		.src31_valid         (cmd_xbar_demux_001_src31_valid),         //          .valid
		.src31_data          (cmd_xbar_demux_001_src31_data),          //          .data
		.src31_channel       (cmd_xbar_demux_001_src31_channel),       //          .channel
		.src31_startofpacket (cmd_xbar_demux_001_src31_startofpacket), //          .startofpacket
		.src31_endofpacket   (cmd_xbar_demux_001_src31_endofpacket),   //          .endofpacket
		.src32_ready         (cmd_xbar_demux_001_src32_ready),         //     src32.ready
		.src32_valid         (cmd_xbar_demux_001_src32_valid),         //          .valid
		.src32_data          (cmd_xbar_demux_001_src32_data),          //          .data
		.src32_channel       (cmd_xbar_demux_001_src32_channel),       //          .channel
		.src32_startofpacket (cmd_xbar_demux_001_src32_startofpacket), //          .startofpacket
		.src32_endofpacket   (cmd_xbar_demux_001_src32_endofpacket),   //          .endofpacket
		.src33_ready         (cmd_xbar_demux_001_src33_ready),         //     src33.ready
		.src33_valid         (cmd_xbar_demux_001_src33_valid),         //          .valid
		.src33_data          (cmd_xbar_demux_001_src33_data),          //          .data
		.src33_channel       (cmd_xbar_demux_001_src33_channel),       //          .channel
		.src33_startofpacket (cmd_xbar_demux_001_src33_startofpacket), //          .startofpacket
		.src33_endofpacket   (cmd_xbar_demux_001_src33_endofpacket),   //          .endofpacket
		.src34_ready         (cmd_xbar_demux_001_src34_ready),         //     src34.ready
		.src34_valid         (cmd_xbar_demux_001_src34_valid),         //          .valid
		.src34_data          (cmd_xbar_demux_001_src34_data),          //          .data
		.src34_channel       (cmd_xbar_demux_001_src34_channel),       //          .channel
		.src34_startofpacket (cmd_xbar_demux_001_src34_startofpacket), //          .startofpacket
		.src34_endofpacket   (cmd_xbar_demux_001_src34_endofpacket),   //          .endofpacket
		.src35_ready         (cmd_xbar_demux_001_src35_ready),         //     src35.ready
		.src35_valid         (cmd_xbar_demux_001_src35_valid),         //          .valid
		.src35_data          (cmd_xbar_demux_001_src35_data),          //          .data
		.src35_channel       (cmd_xbar_demux_001_src35_channel),       //          .channel
		.src35_startofpacket (cmd_xbar_demux_001_src35_startofpacket), //          .startofpacket
		.src35_endofpacket   (cmd_xbar_demux_001_src35_endofpacket),   //          .endofpacket
		.src36_ready         (cmd_xbar_demux_001_src36_ready),         //     src36.ready
		.src36_valid         (cmd_xbar_demux_001_src36_valid),         //          .valid
		.src36_data          (cmd_xbar_demux_001_src36_data),          //          .data
		.src36_channel       (cmd_xbar_demux_001_src36_channel),       //          .channel
		.src36_startofpacket (cmd_xbar_demux_001_src36_startofpacket), //          .startofpacket
		.src36_endofpacket   (cmd_xbar_demux_001_src36_endofpacket),   //          .endofpacket
		.src37_ready         (cmd_xbar_demux_001_src37_ready),         //     src37.ready
		.src37_valid         (cmd_xbar_demux_001_src37_valid),         //          .valid
		.src37_data          (cmd_xbar_demux_001_src37_data),          //          .data
		.src37_channel       (cmd_xbar_demux_001_src37_channel),       //          .channel
		.src37_startofpacket (cmd_xbar_demux_001_src37_startofpacket), //          .startofpacket
		.src37_endofpacket   (cmd_xbar_demux_001_src37_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_004 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (cpu_jtag_debug_module_reset_reset),     // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_005 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (cpu_jtag_debug_module_reset_reset),     // clk_reset.reset
		.sink_ready         (addr_router_005_src_ready),             //      sink.ready
		.sink_channel       (addr_router_005_src_channel),           //          .channel
		.sink_data          (addr_router_005_src_data),              //          .data
		.sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_005_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_006 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_006_src_ready),             //      sink.ready
		.sink_channel       (addr_router_006_src_channel),           //          .channel
		.sink_data          (addr_router_006_src_data),              //          .data
		.sink_startofpacket (addr_router_006_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_006_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_006_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (sys_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (sys_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (sys_clk),                               //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_016 cmd_xbar_mux_016 (
		.clk                 (sys_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_016_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_016_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_016_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_016_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_016_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_016_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_001_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_001_src_valid),           //          .valid
		.sink0_channel       (width_adapter_001_src_channel),         //          .channel
		.sink0_data          (width_adapter_001_src_data),            //          .data
		.sink0_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_004_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (cmd_xbar_demux_005_src0_ready),         //     sink4.ready
		.sink4_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.sink4_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.sink4_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.sink4_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (cmd_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (cmd_xbar_demux_006_src0_ready),         //     sink5.ready
		.sink5_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.sink5_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.sink5_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.sink5_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (cmd_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_006 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_007 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_008 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_009 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_010 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_011 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_012 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_013 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_014 rsp_xbar_demux_014 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_015 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_016 rsp_xbar_demux_016 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_016_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_016_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_016_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_016_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_016_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_016_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_016_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_016_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_016_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_016_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_016_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_016_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_016_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_016_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_016_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_016_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_016_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_016_src3_endofpacket),   //          .endofpacket
		.src4_ready         (rsp_xbar_demux_016_src4_ready),         //      src4.ready
		.src4_valid         (rsp_xbar_demux_016_src4_valid),         //          .valid
		.src4_data          (rsp_xbar_demux_016_src4_data),          //          .data
		.src4_channel       (rsp_xbar_demux_016_src4_channel),       //          .channel
		.src4_startofpacket (rsp_xbar_demux_016_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (rsp_xbar_demux_016_src4_endofpacket),   //          .endofpacket
		.src5_ready         (rsp_xbar_demux_016_src5_ready),         //      src5.ready
		.src5_valid         (rsp_xbar_demux_016_src5_valid),         //          .valid
		.src5_data          (rsp_xbar_demux_016_src5_data),          //          .data
		.src5_channel       (rsp_xbar_demux_016_src5_channel),       //          .channel
		.src5_startofpacket (rsp_xbar_demux_016_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (rsp_xbar_demux_016_src5_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_017 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_014 rsp_xbar_demux_018 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_019 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_020 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_021 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_022 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_023 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_024 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_025 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_026 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_026_src_ready),               //      sink.ready
		.sink_channel       (id_router_026_src_channel),             //          .channel
		.sink_data          (id_router_026_src_data),                //          .data
		.sink_startofpacket (id_router_026_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_026_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_026_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_027 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_027_src_ready),               //      sink.ready
		.sink_channel       (id_router_027_src_channel),             //          .channel
		.sink_data          (id_router_027_src_data),                //          .data
		.sink_startofpacket (id_router_027_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_027_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_027_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_014 rsp_xbar_demux_028 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_028_src_ready),               //      sink.ready
		.sink_channel       (id_router_028_src_channel),             //          .channel
		.sink_data          (id_router_028_src_data),                //          .data
		.sink_startofpacket (id_router_028_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_028_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_028_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_029 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_029_src_ready),               //      sink.ready
		.sink_channel       (id_router_029_src_channel),             //          .channel
		.sink_data          (id_router_029_src_data),                //          .data
		.sink_startofpacket (id_router_029_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_029_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_029_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_029_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_030 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_030_src_ready),               //      sink.ready
		.sink_channel       (id_router_030_src_channel),             //          .channel
		.sink_data          (id_router_030_src_data),                //          .data
		.sink_startofpacket (id_router_030_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_030_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_030_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_030_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_030_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_014 rsp_xbar_demux_031 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_031_src_ready),               //      sink.ready
		.sink_channel       (id_router_031_src_channel),             //          .channel
		.sink_data          (id_router_031_src_data),                //          .data
		.sink_startofpacket (id_router_031_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_031_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_031_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_031_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_031_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_032 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_032_src_ready),               //      sink.ready
		.sink_channel       (id_router_032_src_channel),             //          .channel
		.sink_data          (id_router_032_src_data),                //          .data
		.sink_startofpacket (id_router_032_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_032_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_032_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_032_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_032_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_033 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_033_src_ready),               //      sink.ready
		.sink_channel       (id_router_033_src_channel),             //          .channel
		.sink_data          (id_router_033_src_data),                //          .data
		.sink_startofpacket (id_router_033_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_033_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_033_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_033_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_033_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_034 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_034_src_ready),               //      sink.ready
		.sink_channel       (id_router_034_src_channel),             //          .channel
		.sink_data          (id_router_034_src_data),                //          .data
		.sink_startofpacket (id_router_034_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_034_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_034_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_034_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_034_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_035 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (cpu_jtag_debug_module_reset_reset),     // clk_reset.reset
		.sink_ready         (id_router_035_src_ready),               //      sink.ready
		.sink_channel       (id_router_035_src_channel),             //          .channel
		.sink_data          (id_router_035_src_data),                //          .data
		.sink_startofpacket (id_router_035_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_035_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_035_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_035_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_035_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_036 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (cpu_jtag_debug_module_reset_reset),     // clk_reset.reset
		.sink_ready         (id_router_036_src_ready),               //      sink.ready
		.sink_channel       (id_router_036_src_channel),             //          .channel
		.sink_data          (id_router_036_src_data),                //          .data
		.sink_startofpacket (id_router_036_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_036_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_036_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_036_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_036_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_037 (
		.clk                (sys_clk),                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_037_src_ready),               //      sink.ready
		.sink_channel       (id_router_037_src_channel),             //          .channel
		.sink_data          (id_router_037_src_data),                //          .data
		.sink_startofpacket (id_router_037_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_037_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_037_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_037_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_037_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (sys_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (sys_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (width_adapter_005_src_ready),           //    sink14.ready
		.sink14_valid         (width_adapter_005_src_valid),           //          .valid
		.sink14_channel       (width_adapter_005_src_channel),         //          .channel
		.sink14_data          (width_adapter_005_src_data),            //          .data
		.sink14_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink14_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (width_adapter_006_src_ready),           //    sink16.ready
		.sink16_valid         (width_adapter_006_src_valid),           //          .valid
		.sink16_channel       (width_adapter_006_src_channel),         //          .channel
		.sink16_data          (width_adapter_006_src_data),            //          .data
		.sink16_startofpacket (width_adapter_006_src_startofpacket),   //          .startofpacket
		.sink16_endofpacket   (width_adapter_006_src_endofpacket),     //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (width_adapter_007_src_ready),           //    sink18.ready
		.sink18_valid         (width_adapter_007_src_valid),           //          .valid
		.sink18_channel       (width_adapter_007_src_channel),         //          .channel
		.sink18_data          (width_adapter_007_src_data),            //          .data
		.sink18_startofpacket (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink18_endofpacket   (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_022_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_023_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink24_ready         (rsp_xbar_demux_024_src0_ready),         //    sink24.ready
		.sink24_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink24_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink24_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink24_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink24_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink25_ready         (rsp_xbar_demux_025_src0_ready),         //    sink25.ready
		.sink25_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink25_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink25_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.sink25_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink25_endofpacket   (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.sink26_ready         (rsp_xbar_demux_026_src0_ready),         //    sink26.ready
		.sink26_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.sink26_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.sink26_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.sink26_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.sink26_endofpacket   (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.sink27_ready         (rsp_xbar_demux_027_src0_ready),         //    sink27.ready
		.sink27_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.sink27_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.sink27_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.sink27_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.sink27_endofpacket   (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.sink28_ready         (width_adapter_008_src_ready),           //    sink28.ready
		.sink28_valid         (width_adapter_008_src_valid),           //          .valid
		.sink28_channel       (width_adapter_008_src_channel),         //          .channel
		.sink28_data          (width_adapter_008_src_data),            //          .data
		.sink28_startofpacket (width_adapter_008_src_startofpacket),   //          .startofpacket
		.sink28_endofpacket   (width_adapter_008_src_endofpacket),     //          .endofpacket
		.sink29_ready         (rsp_xbar_demux_029_src0_ready),         //    sink29.ready
		.sink29_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.sink29_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.sink29_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.sink29_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.sink29_endofpacket   (rsp_xbar_demux_029_src0_endofpacket),   //          .endofpacket
		.sink30_ready         (rsp_xbar_demux_030_src0_ready),         //    sink30.ready
		.sink30_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.sink30_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.sink30_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.sink30_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.sink30_endofpacket   (rsp_xbar_demux_030_src0_endofpacket),   //          .endofpacket
		.sink31_ready         (width_adapter_009_src_ready),           //    sink31.ready
		.sink31_valid         (width_adapter_009_src_valid),           //          .valid
		.sink31_channel       (width_adapter_009_src_channel),         //          .channel
		.sink31_data          (width_adapter_009_src_data),            //          .data
		.sink31_startofpacket (width_adapter_009_src_startofpacket),   //          .startofpacket
		.sink31_endofpacket   (width_adapter_009_src_endofpacket),     //          .endofpacket
		.sink32_ready         (rsp_xbar_demux_032_src0_ready),         //    sink32.ready
		.sink32_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.sink32_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.sink32_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.sink32_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.sink32_endofpacket   (rsp_xbar_demux_032_src0_endofpacket),   //          .endofpacket
		.sink33_ready         (rsp_xbar_demux_033_src0_ready),         //    sink33.ready
		.sink33_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.sink33_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.sink33_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.sink33_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.sink33_endofpacket   (rsp_xbar_demux_033_src0_endofpacket),   //          .endofpacket
		.sink34_ready         (rsp_xbar_demux_034_src0_ready),         //    sink34.ready
		.sink34_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.sink34_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.sink34_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.sink34_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.sink34_endofpacket   (rsp_xbar_demux_034_src0_endofpacket),   //          .endofpacket
		.sink35_ready         (rsp_xbar_demux_035_src0_ready),         //    sink35.ready
		.sink35_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.sink35_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.sink35_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.sink35_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.sink35_endofpacket   (rsp_xbar_demux_035_src0_endofpacket),   //          .endofpacket
		.sink36_ready         (rsp_xbar_demux_036_src0_ready),         //    sink36.ready
		.sink36_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.sink36_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.sink36_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.sink36_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.sink36_endofpacket   (rsp_xbar_demux_036_src0_endofpacket),   //          .endofpacket
		.sink37_ready         (rsp_xbar_demux_037_src0_ready),         //    sink37.ready
		.sink37_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.sink37_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.sink37_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.sink37_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.sink37_endofpacket   (rsp_xbar_demux_037_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (110),
		.IN_PKT_RESPONSE_STATUS_L      (109),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (111),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (83),
		.OUT_PKT_RESPONSE_STATUS_L     (82),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (38),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (sys_clk),                                //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src14_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src14_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src14_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src14_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),          //       src.endofpacket
		.out_data             (width_adapter_src_data),                 //          .data
		.out_channel          (width_adapter_src_channel),              //          .channel
		.out_valid            (width_adapter_src_valid),                //          .valid
		.out_ready            (width_adapter_src_ready),                //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),        //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (110),
		.IN_PKT_RESPONSE_STATUS_L      (109),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (111),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (92),
		.OUT_PKT_RESPONSE_STATUS_L     (91),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (38),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_001 (
		.clk                  (sys_clk),                                //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src16_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src16_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src16_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src16_data),          //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_001_src_data),             //          .data
		.out_channel          (width_adapter_001_src_channel),          //          .channel
		.out_valid            (width_adapter_001_src_valid),            //          .valid
		.out_ready            (width_adapter_001_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (110),
		.IN_PKT_RESPONSE_STATUS_L      (109),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (111),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (83),
		.OUT_PKT_RESPONSE_STATUS_L     (82),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (38),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (sys_clk),                                //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src18_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src18_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src18_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src18_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src18_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_002_src_data),             //          .data
		.out_channel          (width_adapter_002_src_channel),          //          .channel
		.out_valid            (width_adapter_002_src_valid),            //          .valid
		.out_ready            (width_adapter_002_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (110),
		.IN_PKT_RESPONSE_STATUS_L      (109),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (111),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (83),
		.OUT_PKT_RESPONSE_STATUS_L     (82),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (38),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_003 (
		.clk                  (sys_clk),                                //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src28_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src28_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src28_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src28_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src28_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src28_data),          //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_003_src_data),             //          .data
		.out_channel          (width_adapter_003_src_channel),          //          .channel
		.out_valid            (width_adapter_003_src_valid),            //          .valid
		.out_ready            (width_adapter_003_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (110),
		.IN_PKT_RESPONSE_STATUS_L      (109),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (111),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (83),
		.OUT_PKT_RESPONSE_STATUS_L     (82),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (38),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_004 (
		.clk                  (sys_clk),                                //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src31_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src31_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src31_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src31_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src31_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src31_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_004_src_data),             //          .data
		.out_channel          (width_adapter_004_src_channel),          //          .channel
		.out_valid            (width_adapter_004_src_valid),            //          .valid
		.out_ready            (width_adapter_004_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (83),
		.IN_PKT_RESPONSE_STATUS_L      (82),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (110),
		.OUT_PKT_RESPONSE_STATUS_L     (109),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (111),
		.ST_CHANNEL_W                  (38),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_005 (
		.clk                  (sys_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_014_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_014_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_014_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_014_src0_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (92),
		.IN_PKT_RESPONSE_STATUS_L      (91),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (110),
		.OUT_PKT_RESPONSE_STATUS_L     (109),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (111),
		.ST_CHANNEL_W                  (38),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_006 (
		.clk                  (sys_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_016_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_016_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_016_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_016_src0_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_006_src_data),            //          .data
		.out_channel          (width_adapter_006_src_channel),         //          .channel
		.out_valid            (width_adapter_006_src_valid),           //          .valid
		.out_ready            (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (83),
		.IN_PKT_RESPONSE_STATUS_L      (82),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (110),
		.OUT_PKT_RESPONSE_STATUS_L     (109),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (111),
		.ST_CHANNEL_W                  (38),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_007 (
		.clk                  (sys_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_018_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_018_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_018_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_018_src0_data),          //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_007_src_data),            //          .data
		.out_channel          (width_adapter_007_src_channel),         //          .channel
		.out_valid            (width_adapter_007_src_valid),           //          .valid
		.out_ready            (width_adapter_007_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (83),
		.IN_PKT_RESPONSE_STATUS_L      (82),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (110),
		.OUT_PKT_RESPONSE_STATUS_L     (109),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (111),
		.ST_CHANNEL_W                  (38),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_008 (
		.clk                  (sys_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_028_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_028_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_028_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_028_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_028_src0_data),          //          .data
		.out_endofpacket      (width_adapter_008_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_008_src_data),            //          .data
		.out_channel          (width_adapter_008_src_channel),         //          .channel
		.out_valid            (width_adapter_008_src_valid),           //          .valid
		.out_ready            (width_adapter_008_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_008_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (83),
		.IN_PKT_RESPONSE_STATUS_L      (82),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (110),
		.OUT_PKT_RESPONSE_STATUS_L     (109),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (111),
		.ST_CHANNEL_W                  (38),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_009 (
		.clk                  (sys_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_031_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_031_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_031_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_031_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_031_src0_data),          //          .data
		.out_endofpacket      (width_adapter_009_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_009_src_data),            //          .data
		.out_channel          (width_adapter_009_src_channel),         //          .channel
		.out_valid            (width_adapter_009_src_valid),           //          .valid
		.out_ready            (width_adapter_009_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_009_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	nios_system_irq_mapper irq_mapper (
		.clk            (sys_clk),                        //        clk.clk
		.reset          (rst_controller_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),       //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),       //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),       //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),       //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),       //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),       //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),       //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),       //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),       //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),       //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),      // receiver10.irq
		.receiver11_irq (irq_mapper_receiver11_irq),      // receiver11.irq
		.sender_irq     (cpu_d_irq_irq)                   //     sender.irq
	);

	nios_system_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (2),
		.outErrorWidth   (6),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (sys_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_005_reset_out_reset),    // in_rst_0.reset
		.in_0_ready          (enet_receive_ready),                    //     in_0.ready
		.in_0_valid          (enet_receive_valid),                    //         .valid
		.in_0_data           (enet_receive_data),                     //         .data
		.in_0_startofpacket  (enet_receive_startofpacket),            //         .startofpacket
		.in_0_endofpacket    (enet_receive_endofpacket),              //         .endofpacket
		.in_0_empty          (enet_receive_empty),                    //         .empty
		.in_0_error          (enet_receive_error),                    //         .error
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //    out_0.ready
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_data          (avalon_st_adapter_out_0_data),          //         .data
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_channel       (avalon_st_adapter_out_0_channel),       //         .channel
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	nios_system_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (2),
		.inErrorWidth    (6),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (sys_clk),                                                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_006_reset_out_reset),                            // in_rst_0.reset
		.in_0_ready          (videoconferencing_dma_0_avalon_streaming_source_ready),         //     in_0.ready
		.in_0_valid          (videoconferencing_dma_0_avalon_streaming_source_valid),         //         .valid
		.in_0_data           (videoconferencing_dma_0_avalon_streaming_source_data),          //         .data
		.in_0_startofpacket  (videoconferencing_dma_0_avalon_streaming_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (videoconferencing_dma_0_avalon_streaming_source_endofpacket),   //         .endofpacket
		.in_0_channel        (videoconferencing_dma_0_avalon_streaming_source_channel),       //         .channel
		.in_0_error          (videoconferencing_dma_0_avalon_streaming_source_error),         //         .error
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),                             //    out_0.ready
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),                             //         .valid
		.out_0_data          (avalon_st_adapter_001_out_0_data),                              //         .data
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket),                     //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),                       //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty),                             //         .empty
		.out_0_error         (avalon_st_adapter_001_out_0_error)                              //         .error
	);

endmodule
