// nios_system_tb.v

// Generated using ACDS version 13.0sp1 232 at 2015.05.15.21:27:45

`timescale 1 ps / 1 ps
module nios_system_tb (
	);

	wire         nios_system_inst_clk_clk_in_bfm_clk_clk;                                // nios_system_inst_clk_clk_in_bfm:clk -> [nios_system_inst:clk, nios_system_inst_merged_resets_in_reset_bfm:clk]
	wire         nios_system_inst_clk_27_clk_in_bfm_clk_clk;                             // nios_system_inst_clk_27_clk_in_bfm:clk -> nios_system_inst:clk_27
	wire         nios_system_inst_enet_pcs_mac_tx_bfm_clk_clk;                           // nios_system_inst_enet_pcs_mac_tx_bfm:clk -> nios_system_inst:enet_pcs_mac_tx_clk
	wire         nios_system_inst_enet_pcs_mac_rx_bfm_clk_clk;                           // nios_system_inst_enet_pcs_mac_rx_bfm:clk -> nios_system_inst:enet_pcs_mac_rx_clk
	wire         nios_system_inst_merged_resets_in_reset_bfm_reset_reset;                // nios_system_inst_merged_resets_in_reset_bfm:reset -> nios_system_inst:reset_n
	wire   [6:0] nios_system_inst_hex7_hex4_external_interface_hex6;                     // nios_system_inst:HEX6_from_the_HEX7_HEX4 -> nios_system_inst_HEX7_HEX4_external_interface_bfm:sig_HEX6
	wire   [6:0] nios_system_inst_hex7_hex4_external_interface_hex5;                     // nios_system_inst:HEX5_from_the_HEX7_HEX4 -> nios_system_inst_HEX7_HEX4_external_interface_bfm:sig_HEX5
	wire   [6:0] nios_system_inst_hex7_hex4_external_interface_hex4;                     // nios_system_inst:HEX4_from_the_HEX7_HEX4 -> nios_system_inst_HEX7_HEX4_external_interface_bfm:sig_HEX4
	wire   [6:0] nios_system_inst_hex7_hex4_external_interface_hex7;                     // nios_system_inst:HEX7_from_the_HEX7_HEX4 -> nios_system_inst_HEX7_HEX4_external_interface_bfm:sig_HEX7
	wire  [15:0] nios_system_inst_sram_external_interface_dq;                            // [] -> [nios_system_inst:SRAM_DQ_to_and_from_the_SRAM, nios_system_inst_SRAM_external_interface_bfm:sig_DQ]
	wire         nios_system_inst_sram_external_interface_ce_n;                          // nios_system_inst:SRAM_CE_N_from_the_SRAM -> nios_system_inst_SRAM_external_interface_bfm:sig_CE_N
	wire         nios_system_inst_sram_external_interface_ub_n;                          // nios_system_inst:SRAM_UB_N_from_the_SRAM -> nios_system_inst_SRAM_external_interface_bfm:sig_UB_N
	wire         nios_system_inst_sram_external_interface_oe_n;                          // nios_system_inst:SRAM_OE_N_from_the_SRAM -> nios_system_inst_SRAM_external_interface_bfm:sig_OE_N
	wire         nios_system_inst_sram_external_interface_lb_n;                          // nios_system_inst:SRAM_LB_N_from_the_SRAM -> nios_system_inst_SRAM_external_interface_bfm:sig_LB_N
	wire         nios_system_inst_sram_external_interface_we_n;                          // nios_system_inst:SRAM_WE_N_from_the_SRAM -> nios_system_inst_SRAM_external_interface_bfm:sig_WE_N
	wire  [19:0] nios_system_inst_sram_external_interface_addr;                          // nios_system_inst:SRAM_ADDR_from_the_SRAM -> nios_system_inst_SRAM_external_interface_bfm:sig_ADDR
	wire         nios_system_inst_char_lcd_16x2_external_interface_rs;                   // nios_system_inst:LCD_RS_from_the_Char_LCD_16x2 -> nios_system_inst_Char_LCD_16x2_external_interface_bfm:sig_RS
	wire         nios_system_inst_char_lcd_16x2_external_interface_on;                   // nios_system_inst:LCD_ON_from_the_Char_LCD_16x2 -> nios_system_inst_Char_LCD_16x2_external_interface_bfm:sig_ON
	wire         nios_system_inst_char_lcd_16x2_external_interface_en;                   // nios_system_inst:LCD_EN_from_the_Char_LCD_16x2 -> nios_system_inst_Char_LCD_16x2_external_interface_bfm:sig_EN
	wire         nios_system_inst_char_lcd_16x2_external_interface_blon;                 // nios_system_inst:LCD_BLON_from_the_Char_LCD_16x2 -> nios_system_inst_Char_LCD_16x2_external_interface_bfm:sig_BLON
	wire         nios_system_inst_char_lcd_16x2_external_interface_rw;                   // nios_system_inst:LCD_RW_from_the_Char_LCD_16x2 -> nios_system_inst_Char_LCD_16x2_external_interface_bfm:sig_RW
	wire   [7:0] nios_system_inst_char_lcd_16x2_external_interface_data;                 // [] -> [nios_system_inst:LCD_DATA_to_and_from_the_Char_LCD_16x2, nios_system_inst_Char_LCD_16x2_external_interface_bfm:sig_DATA]
	wire         nios_system_inst_serial_port_external_interface_bfm_conduit_rxd;        // nios_system_inst_Serial_Port_external_interface_bfm:sig_RXD -> nios_system_inst:UART_RXD_to_the_Serial_Port
	wire         nios_system_inst_serial_port_external_interface_txd;                    // nios_system_inst:UART_TXD_from_the_Serial_Port -> nios_system_inst_Serial_Port_external_interface_bfm:sig_TXD
	wire         nios_system_inst_audio_external_interface_bfm_conduit_adclrck;          // nios_system_inst_Audio_external_interface_bfm:sig_ADCLRCK -> nios_system_inst:AUD_ADCLRCK_to_the_Audio
	wire         nios_system_inst_audio_external_interface_bfm_conduit_adcdat;           // nios_system_inst_Audio_external_interface_bfm:sig_ADCDAT -> nios_system_inst:AUD_ADCDAT_to_the_Audio
	wire         nios_system_inst_audio_external_interface_bfm_conduit_daclrck;          // nios_system_inst_Audio_external_interface_bfm:sig_DACLRCK -> nios_system_inst:AUD_DACLRCK_to_the_Audio
	wire         nios_system_inst_audio_external_interface_dacdat;                       // nios_system_inst:AUD_DACDAT_from_the_Audio -> nios_system_inst_Audio_external_interface_bfm:sig_DACDAT
	wire         nios_system_inst_audio_external_interface_bfm_conduit_bclk;             // nios_system_inst_Audio_external_interface_bfm:sig_BCLK -> nios_system_inst:AUD_BCLK_to_the_Audio
	wire  [17:0] nios_system_inst_red_leds_external_interface_export;                    // nios_system_inst:LEDR_from_the_Red_LEDs -> nios_system_inst_Red_LEDs_external_interface_bfm:sig_export
	wire         nios_system_inst_sdram_wire_cs_n;                                       // nios_system_inst:zs_cs_n_from_the_SDRAM -> nios_system_inst_SDRAM_wire_bfm:sig_cs_n
	wire   [1:0] nios_system_inst_sdram_wire_ba;                                         // nios_system_inst:zs_ba_from_the_SDRAM -> nios_system_inst_SDRAM_wire_bfm:sig_ba
	wire   [3:0] nios_system_inst_sdram_wire_dqm;                                        // nios_system_inst:zs_dqm_from_the_SDRAM -> nios_system_inst_SDRAM_wire_bfm:sig_dqm
	wire         nios_system_inst_sdram_wire_cke;                                        // nios_system_inst:zs_cke_from_the_SDRAM -> nios_system_inst_SDRAM_wire_bfm:sig_cke
	wire  [12:0] nios_system_inst_sdram_wire_addr;                                       // nios_system_inst:zs_addr_from_the_SDRAM -> nios_system_inst_SDRAM_wire_bfm:sig_addr
	wire         nios_system_inst_sdram_wire_we_n;                                       // nios_system_inst:zs_we_n_from_the_SDRAM -> nios_system_inst_SDRAM_wire_bfm:sig_we_n
	wire         nios_system_inst_sdram_wire_ras_n;                                      // nios_system_inst:zs_ras_n_from_the_SDRAM -> nios_system_inst_SDRAM_wire_bfm:sig_ras_n
	wire  [31:0] nios_system_inst_sdram_wire_dq;                                         // [] -> [nios_system_inst:zs_dq_to_and_from_the_SDRAM, nios_system_inst_SDRAM_wire_bfm:sig_dq]
	wire         nios_system_inst_sdram_wire_cas_n;                                      // nios_system_inst:zs_cas_n_from_the_SDRAM -> nios_system_inst_SDRAM_wire_bfm:sig_cas_n
	wire  [31:0] nios_system_inst_expansion_jp5_external_interface_export;               // [] -> [nios_system_inst:GPIO_to_and_from_the_Expansion_JP5, nios_system_inst_Expansion_JP5_external_interface_bfm:sig_export]
	wire   [8:0] nios_system_inst_green_leds_external_interface_export;                  // nios_system_inst:LEDG_from_the_Green_LEDs -> nios_system_inst_Green_LEDs_external_interface_bfm:sig_export
	wire         nios_system_inst_ps2_port_dual_external_interface_clk;                  // [] -> [nios_system_inst:PS2_CLK_to_and_from_the_PS2_Port_Dual, nios_system_inst_PS2_Port_Dual_external_interface_bfm:sig_CLK]
	wire         nios_system_inst_ps2_port_dual_external_interface_dat;                  // [] -> [nios_system_inst:PS2_DAT_to_and_from_the_PS2_Port_Dual, nios_system_inst_PS2_Port_Dual_external_interface_bfm:sig_DAT]
	wire  [17:0] nios_system_inst_slider_switches_external_interface_bfm_conduit_export; // nios_system_inst_Slider_Switches_external_interface_bfm:sig_export -> nios_system_inst:Slider_Switches_external_interface_export
	wire         nios_system_inst_av_config_external_interface_sclk;                     // nios_system_inst:I2C_SCLK_from_the_AV_Config -> nios_system_inst_AV_Config_external_interface_bfm:sig_SCLK
	wire         nios_system_inst_av_config_external_interface_sdat;                     // [] -> [nios_system_inst:I2C_SDAT_to_and_from_the_AV_Config, nios_system_inst_AV_Config_external_interface_bfm:sig_SDAT]
	wire         nios_system_inst_ps2_port_external_interface_clk;                       // [] -> [nios_system_inst:PS2_CLK_to_and_from_the_PS2_Port, nios_system_inst_PS2_Port_external_interface_bfm:sig_CLK]
	wire         nios_system_inst_ps2_port_external_interface_dat;                       // [] -> [nios_system_inst:PS2_DAT_to_and_from_the_PS2_Port, nios_system_inst_PS2_Port_external_interface_bfm:sig_DAT]
	wire   [3:0] nios_system_inst_pushbuttons_external_interface_bfm_conduit_export;     // nios_system_inst_Pushbuttons_external_interface_bfm:sig_export -> nios_system_inst:KEY_to_the_Pushbuttons
	wire   [6:0] nios_system_inst_hex3_hex0_external_interface_hex2;                     // nios_system_inst:HEX2_from_the_HEX3_HEX0 -> nios_system_inst_HEX3_HEX0_external_interface_bfm:sig_HEX2
	wire   [6:0] nios_system_inst_hex3_hex0_external_interface_hex1;                     // nios_system_inst:HEX1_from_the_HEX3_HEX0 -> nios_system_inst_HEX3_HEX0_external_interface_bfm:sig_HEX1
	wire   [6:0] nios_system_inst_hex3_hex0_external_interface_hex0;                     // nios_system_inst:HEX0_from_the_HEX3_HEX0 -> nios_system_inst_HEX3_HEX0_external_interface_bfm:sig_HEX0
	wire   [6:0] nios_system_inst_hex3_hex0_external_interface_hex3;                     // nios_system_inst:HEX3_from_the_HEX3_HEX0 -> nios_system_inst_HEX3_HEX0_external_interface_bfm:sig_HEX3
	wire         nios_system_inst_irda_bfm_conduit_rxd;                                  // nios_system_inst_irda_bfm:sig_RXD -> nios_system_inst:irda_RXD
	wire         nios_system_inst_irda_txd;                                              // nios_system_inst:irda_TXD -> nios_system_inst_irda_bfm:sig_TXD
	wire         nios_system_inst_sdcard_b_sd_dat;                                       // [] -> [nios_system_inst:sdcard_b_SD_dat, nios_system_inst_sdcard_bfm:sig_b_SD_dat]
	wire         nios_system_inst_sdcard_b_sd_cmd;                                       // [] -> [nios_system_inst:sdcard_b_SD_cmd, nios_system_inst_sdcard_bfm:sig_b_SD_cmd]
	wire         nios_system_inst_sdcard_o_sd_clock;                                     // nios_system_inst:sdcard_o_SD_clock -> nios_system_inst_sdcard_bfm:sig_o_SD_clock
	wire         nios_system_inst_sdcard_b_sd_dat3;                                      // [] -> [nios_system_inst:sdcard_b_SD_dat3, nios_system_inst_sdcard_bfm:sig_b_SD_dat3]
	wire   [7:0] nios_system_inst_flash_dq;                                              // [] -> [nios_system_inst:flash_DQ, nios_system_inst_flash_bfm:sig_DQ]
	wire         nios_system_inst_flash_ce_n;                                            // nios_system_inst:flash_CE_N -> nios_system_inst_flash_bfm:sig_CE_N
	wire         nios_system_inst_flash_oe_n;                                            // nios_system_inst:flash_OE_N -> nios_system_inst_flash_bfm:sig_OE_N
	wire         nios_system_inst_flash_we_n;                                            // nios_system_inst:flash_WE_N -> nios_system_inst_flash_bfm:sig_WE_N
	wire  [22:0] nios_system_inst_flash_addr;                                            // nios_system_inst:flash_ADDR -> nios_system_inst_flash_bfm:sig_ADDR
	wire         nios_system_inst_flash_rst_n;                                           // nios_system_inst:flash_RST_N -> nios_system_inst_flash_bfm:sig_RST_N
	wire         nios_system_inst_video_in_bfm_conduit_td_clk27;                         // nios_system_inst_video_in_bfm:sig_TD_CLK27 -> nios_system_inst:video_in_TD_CLK27
	wire         nios_system_inst_video_in_bfm_conduit_td_hs;                            // nios_system_inst_video_in_bfm:sig_TD_HS -> nios_system_inst:video_in_TD_HS
	wire         nios_system_inst_video_in_td_reset;                                     // nios_system_inst:video_in_TD_RESET -> nios_system_inst_video_in_bfm:sig_TD_RESET
	wire         nios_system_inst_video_in_bfm_conduit_clk27_reset;                      // nios_system_inst_video_in_bfm:sig_clk27_reset -> nios_system_inst:video_in_clk27_reset
	wire   [7:0] nios_system_inst_video_in_bfm_conduit_td_data;                          // nios_system_inst_video_in_bfm:sig_TD_DATA -> nios_system_inst:video_in_TD_DATA
	wire         nios_system_inst_video_in_overflow_flag;                                // nios_system_inst:video_in_overflow_flag -> nios_system_inst_video_in_bfm:sig_overflow_flag
	wire         nios_system_inst_video_in_bfm_conduit_td_vs;                            // nios_system_inst_video_in_bfm:sig_TD_VS -> nios_system_inst:video_in_TD_VS
	wire  [15:0] nios_system_inst_camera_config_bfm_conduit_exposure;                    // nios_system_inst_camera_config_bfm:sig_exposure -> nios_system_inst:camera_config_exposure
	wire         nios_system_inst_camera_config_i2c_sdat;                                // [] -> [nios_system_inst:camera_config_I2C_SDAT, nios_system_inst_camera_config_bfm:sig_I2C_SDAT]
	wire         nios_system_inst_camera_config_i2c_sclk;                                // nios_system_inst:camera_config_I2C_SCLK -> nios_system_inst_camera_config_bfm:sig_I2C_SCLK
	wire         nios_system_inst_camera_in_bfm_conduit_line_valid;                      // nios_system_inst_camera_in_bfm:sig_LINE_VALID -> nios_system_inst:camera_in_LINE_VALID
	wire         nios_system_inst_camera_in_bfm_conduit_pixel_clk_reset;                 // nios_system_inst_camera_in_bfm:sig_pixel_clk_reset -> nios_system_inst:camera_in_pixel_clk_reset
	wire         nios_system_inst_camera_in_bfm_conduit_frame_valid;                     // nios_system_inst_camera_in_bfm:sig_FRAME_VALID -> nios_system_inst:camera_in_FRAME_VALID
	wire  [11:0] nios_system_inst_camera_in_bfm_conduit_pixel_data;                      // nios_system_inst_camera_in_bfm:sig_PIXEL_DATA -> nios_system_inst:camera_in_PIXEL_DATA
	wire         nios_system_inst_camera_in_bfm_conduit_pixel_clk;                       // nios_system_inst_camera_in_bfm:sig_PIXEL_CLK -> nios_system_inst:camera_in_PIXEL_CLK
	wire         nios_system_inst_lcd_controller_external_interface_data_en;             // nios_system_inst:lcd_controller_external_interface_DATA_EN -> nios_system_inst_lcd_controller_external_interface_bfm:sig_DATA_EN
	wire   [7:0] nios_system_inst_lcd_controller_external_interface_g;                   // nios_system_inst:lcd_controller_external_interface_G -> nios_system_inst_lcd_controller_external_interface_bfm:sig_G
	wire         nios_system_inst_lcd_controller_external_interface_vs;                  // nios_system_inst:lcd_controller_external_interface_VS -> nios_system_inst_lcd_controller_external_interface_bfm:sig_VS
	wire   [7:0] nios_system_inst_lcd_controller_external_interface_b;                   // nios_system_inst:lcd_controller_external_interface_B -> nios_system_inst_lcd_controller_external_interface_bfm:sig_B
	wire   [7:0] nios_system_inst_lcd_controller_external_interface_r;                   // nios_system_inst:lcd_controller_external_interface_R -> nios_system_inst_lcd_controller_external_interface_bfm:sig_R
	wire         nios_system_inst_lcd_controller_external_interface_hs;                  // nios_system_inst:lcd_controller_external_interface_HS -> nios_system_inst_lcd_controller_external_interface_bfm:sig_HS
	wire         nios_system_inst_lcd_controller_external_interface_clk;                 // nios_system_inst:lcd_controller_external_interface_CLK -> nios_system_inst_lcd_controller_external_interface_bfm:sig_CLK
	wire         nios_system_inst_accelerometer_i2c_sdat;                                // [] -> [nios_system_inst:accelerometer_I2C_SDAT, nios_system_inst_accelerometer_bfm:sig_I2C_SDAT]
	wire         nios_system_inst_accelerometer_bfm_conduit_g_sensor_int;                // nios_system_inst_accelerometer_bfm:sig_G_SENSOR_INT -> nios_system_inst:accelerometer_G_SENSOR_INT
	wire         nios_system_inst_accelerometer_i2c_sclk;                                // nios_system_inst:accelerometer_I2C_SCLK -> nios_system_inst_accelerometer_bfm:sig_I2C_SCLK
	wire         nios_system_inst_accelerometer_g_sensor_cs_n;                           // nios_system_inst:accelerometer_G_SENSOR_CS_N -> nios_system_inst_accelerometer_bfm:sig_G_SENSOR_CS_N
	wire         nios_system_inst_usb_wr_n;                                              // nios_system_inst:usb_WR_N -> nios_system_inst_usb_bfm:sig_WR_N
	wire         nios_system_inst_usb_bfm_conduit_int0;                                  // nios_system_inst_usb_bfm:sig_INT0 -> nios_system_inst:usb_INT0
	wire         nios_system_inst_usb_cs_n;                                              // nios_system_inst:usb_CS_N -> nios_system_inst_usb_bfm:sig_CS_N
	wire         nios_system_inst_usb_bfm_conduit_int1;                                  // nios_system_inst_usb_bfm:sig_INT1 -> nios_system_inst:usb_INT1
	wire   [1:0] nios_system_inst_usb_addr;                                              // nios_system_inst:usb_ADDR -> nios_system_inst_usb_bfm:sig_ADDR
	wire  [15:0] nios_system_inst_usb_data;                                              // [] -> [nios_system_inst:usb_DATA, nios_system_inst_usb_bfm:sig_DATA]
	wire         nios_system_inst_usb_rst_n;                                             // nios_system_inst:usb_RST_N -> nios_system_inst_usb_bfm:sig_RST_N
	wire         nios_system_inst_usb_rd_n;                                              // nios_system_inst:usb_RD_N -> nios_system_inst_usb_bfm:sig_RD_N
	wire   [7:0] nios_system_inst_vga_controller_external_interface_g;                   // nios_system_inst:vga_controller_external_interface_G -> nios_system_inst_vga_controller_external_interface_bfm:sig_G
	wire         nios_system_inst_vga_controller_external_interface_vs;                  // nios_system_inst:vga_controller_external_interface_VS -> nios_system_inst_vga_controller_external_interface_bfm:sig_VS
	wire   [7:0] nios_system_inst_vga_controller_external_interface_b;                   // nios_system_inst:vga_controller_external_interface_B -> nios_system_inst_vga_controller_external_interface_bfm:sig_B
	wire   [7:0] nios_system_inst_vga_controller_external_interface_r;                   // nios_system_inst:vga_controller_external_interface_R -> nios_system_inst_vga_controller_external_interface_bfm:sig_R
	wire         nios_system_inst_vga_controller_external_interface_sync;                // nios_system_inst:vga_controller_external_interface_SYNC -> nios_system_inst_vga_controller_external_interface_bfm:sig_SYNC
	wire         nios_system_inst_vga_controller_external_interface_hs;                  // nios_system_inst:vga_controller_external_interface_HS -> nios_system_inst_vga_controller_external_interface_bfm:sig_HS
	wire         nios_system_inst_vga_controller_external_interface_clk;                 // nios_system_inst:vga_controller_external_interface_CLK -> nios_system_inst_vga_controller_external_interface_bfm:sig_CLK
	wire         nios_system_inst_vga_controller_external_interface_blank;               // nios_system_inst:vga_controller_external_interface_BLANK -> nios_system_inst_vga_controller_external_interface_bfm:sig_BLANK
	wire         nios_system_inst_enet_mac_status_bfm_conduit_set_10;                    // nios_system_inst_enet_mac_status_bfm:sig_set_10 -> nios_system_inst:enet_mac_status_set_10
	wire         nios_system_inst_enet_mac_status_ena_10;                                // nios_system_inst:enet_mac_status_ena_10 -> nios_system_inst_enet_mac_status_bfm:sig_ena_10
	wire         nios_system_inst_enet_mac_status_eth_mode;                              // nios_system_inst:enet_mac_status_eth_mode -> nios_system_inst_enet_mac_status_bfm:sig_eth_mode
	wire         nios_system_inst_enet_mac_status_bfm_conduit_set_1000;                  // nios_system_inst_enet_mac_status_bfm:sig_set_1000 -> nios_system_inst:enet_mac_status_set_1000
	wire   [3:0] nios_system_inst_enet_mac_rgmii_bfm_conduit_rgmii_in;                   // nios_system_inst_enet_mac_rgmii_bfm:sig_rgmii_in -> nios_system_inst:enet_mac_rgmii_rgmii_in
	wire         nios_system_inst_enet_mac_rgmii_tx_control;                             // nios_system_inst:enet_mac_rgmii_tx_control -> nios_system_inst_enet_mac_rgmii_bfm:sig_tx_control
	wire   [3:0] nios_system_inst_enet_mac_rgmii_rgmii_out;                              // nios_system_inst:enet_mac_rgmii_rgmii_out -> nios_system_inst_enet_mac_rgmii_bfm:sig_rgmii_out
	wire         nios_system_inst_enet_mac_rgmii_bfm_conduit_rx_control;                 // nios_system_inst_enet_mac_rgmii_bfm:sig_rx_control -> nios_system_inst:enet_mac_rgmii_rx_control
	wire         nios_system_inst_enet_mac_mdio_bfm_conduit_mdio_in;                     // nios_system_inst_enet_mac_mdio_bfm:sig_mdio_in -> nios_system_inst:enet_mac_mdio_mdio_in
	wire         nios_system_inst_enet_mac_mdio_mdc;                                     // nios_system_inst:enet_mac_mdio_mdc -> nios_system_inst_enet_mac_mdio_bfm:sig_mdc
	wire         nios_system_inst_enet_mac_mdio_mdio_out;                                // nios_system_inst:enet_mac_mdio_mdio_out -> nios_system_inst_enet_mac_mdio_bfm:sig_mdio_out
	wire         nios_system_inst_enet_mac_mdio_mdio_oen;                                // nios_system_inst:enet_mac_mdio_mdio_oen -> nios_system_inst_enet_mac_mdio_bfm:sig_mdio_oen
	wire         nios_system_inst_enet_mac_misc_ff_tx_septy;                             // nios_system_inst:enet_mac_misc_ff_tx_septy -> nios_system_inst_enet_mac_misc_bfm:sig_ff_tx_septy
	wire         nios_system_inst_enet_mac_misc_ff_rx_a_empty;                           // nios_system_inst:enet_mac_misc_ff_rx_a_empty -> nios_system_inst_enet_mac_misc_bfm:sig_ff_rx_a_empty
	wire         nios_system_inst_enet_mac_misc_bfm_conduit_xon_gen;                     // nios_system_inst_enet_mac_misc_bfm:sig_xon_gen -> nios_system_inst:enet_mac_misc_xon_gen
	wire         nios_system_inst_enet_mac_misc_magic_wakeup;                            // nios_system_inst:enet_mac_misc_magic_wakeup -> nios_system_inst_enet_mac_misc_bfm:sig_magic_wakeup
	wire         nios_system_inst_enet_mac_misc_ff_tx_a_full;                            // nios_system_inst:enet_mac_misc_ff_tx_a_full -> nios_system_inst_enet_mac_misc_bfm:sig_ff_tx_a_full
	wire         nios_system_inst_enet_mac_misc_bfm_conduit_xoff_gen;                    // nios_system_inst_enet_mac_misc_bfm:sig_xoff_gen -> nios_system_inst:enet_mac_misc_xoff_gen
	wire         nios_system_inst_enet_mac_misc_bfm_conduit_magic_sleep_n;               // nios_system_inst_enet_mac_misc_bfm:sig_magic_sleep_n -> nios_system_inst:enet_mac_misc_magic_sleep_n
	wire         nios_system_inst_enet_mac_misc_bfm_conduit_ff_tx_crc_fwd;               // nios_system_inst_enet_mac_misc_bfm:sig_ff_tx_crc_fwd -> nios_system_inst:enet_mac_misc_ff_tx_crc_fwd
	wire  [17:0] nios_system_inst_enet_mac_misc_rx_err_stat;                             // nios_system_inst:enet_mac_misc_rx_err_stat -> nios_system_inst_enet_mac_misc_bfm:sig_rx_err_stat
	wire         nios_system_inst_enet_mac_misc_tx_ff_uflow;                             // nios_system_inst:enet_mac_misc_tx_ff_uflow -> nios_system_inst_enet_mac_misc_bfm:sig_tx_ff_uflow
	wire         nios_system_inst_enet_mac_misc_ff_rx_dsav;                              // nios_system_inst:enet_mac_misc_ff_rx_dsav -> nios_system_inst_enet_mac_misc_bfm:sig_ff_rx_dsav
	wire   [3:0] nios_system_inst_enet_mac_misc_rx_frm_type;                             // nios_system_inst:enet_mac_misc_rx_frm_type -> nios_system_inst_enet_mac_misc_bfm:sig_rx_frm_type
	wire         nios_system_inst_enet_mac_misc_ff_rx_a_full;                            // nios_system_inst:enet_mac_misc_ff_rx_a_full -> nios_system_inst_enet_mac_misc_bfm:sig_ff_rx_a_full
	wire         nios_system_inst_enet_mac_misc_ff_tx_a_empty;                           // nios_system_inst:enet_mac_misc_ff_tx_a_empty -> nios_system_inst_enet_mac_misc_bfm:sig_ff_tx_a_empty

	nios_system nios_system_inst (
		.HEX4_from_the_HEX7_HEX4                   (nios_system_inst_hex7_hex4_external_interface_hex4),                     //       HEX7_HEX4_external_interface.HEX4
		.HEX5_from_the_HEX7_HEX4                   (nios_system_inst_hex7_hex4_external_interface_hex5),                     //                                   .HEX5
		.HEX6_from_the_HEX7_HEX4                   (nios_system_inst_hex7_hex4_external_interface_hex6),                     //                                   .HEX6
		.HEX7_from_the_HEX7_HEX4                   (nios_system_inst_hex7_hex4_external_interface_hex7),                     //                                   .HEX7
		.SRAM_DQ_to_and_from_the_SRAM              (nios_system_inst_sram_external_interface_dq),                            //            SRAM_external_interface.DQ
		.SRAM_ADDR_from_the_SRAM                   (nios_system_inst_sram_external_interface_addr),                          //                                   .ADDR
		.SRAM_LB_N_from_the_SRAM                   (nios_system_inst_sram_external_interface_lb_n),                          //                                   .LB_N
		.SRAM_UB_N_from_the_SRAM                   (nios_system_inst_sram_external_interface_ub_n),                          //                                   .UB_N
		.SRAM_CE_N_from_the_SRAM                   (nios_system_inst_sram_external_interface_ce_n),                          //                                   .CE_N
		.SRAM_OE_N_from_the_SRAM                   (nios_system_inst_sram_external_interface_oe_n),                          //                                   .OE_N
		.SRAM_WE_N_from_the_SRAM                   (nios_system_inst_sram_external_interface_we_n),                          //                                   .WE_N
		.LCD_DATA_to_and_from_the_Char_LCD_16x2    (nios_system_inst_char_lcd_16x2_external_interface_data),                 //   Char_LCD_16x2_external_interface.DATA
		.LCD_ON_from_the_Char_LCD_16x2             (nios_system_inst_char_lcd_16x2_external_interface_on),                   //                                   .ON
		.LCD_BLON_from_the_Char_LCD_16x2           (nios_system_inst_char_lcd_16x2_external_interface_blon),                 //                                   .BLON
		.LCD_EN_from_the_Char_LCD_16x2             (nios_system_inst_char_lcd_16x2_external_interface_en),                   //                                   .EN
		.LCD_RS_from_the_Char_LCD_16x2             (nios_system_inst_char_lcd_16x2_external_interface_rs),                   //                                   .RS
		.LCD_RW_from_the_Char_LCD_16x2             (nios_system_inst_char_lcd_16x2_external_interface_rw),                   //                                   .RW
		.sys_clk                                   (),                                                                       //                    sys_clk_out_clk.clk
		.UART_RXD_to_the_Serial_Port               (nios_system_inst_serial_port_external_interface_bfm_conduit_rxd),        //     Serial_Port_external_interface.RXD
		.UART_TXD_from_the_Serial_Port             (nios_system_inst_serial_port_external_interface_txd),                    //                                   .TXD
		.AUD_ADCDAT_to_the_Audio                   (nios_system_inst_audio_external_interface_bfm_conduit_adcdat),           //           Audio_external_interface.ADCDAT
		.AUD_ADCLRCK_to_the_Audio                  (nios_system_inst_audio_external_interface_bfm_conduit_adclrck),          //                                   .ADCLRCK
		.AUD_BCLK_to_the_Audio                     (nios_system_inst_audio_external_interface_bfm_conduit_bclk),             //                                   .BCLK
		.AUD_DACDAT_from_the_Audio                 (nios_system_inst_audio_external_interface_dacdat),                       //                                   .DACDAT
		.AUD_DACLRCK_to_the_Audio                  (nios_system_inst_audio_external_interface_bfm_conduit_daclrck),          //                                   .DACLRCK
		.LEDR_from_the_Red_LEDs                    (nios_system_inst_red_leds_external_interface_export),                    //        Red_LEDs_external_interface.export
		.reset_n                                   (nios_system_inst_merged_resets_in_reset_bfm_reset_reset),                //             merged_resets_in_reset.reset_n
		.zs_addr_from_the_SDRAM                    (nios_system_inst_sdram_wire_addr),                                       //                         SDRAM_wire.addr
		.zs_ba_from_the_SDRAM                      (nios_system_inst_sdram_wire_ba),                                         //                                   .ba
		.zs_cas_n_from_the_SDRAM                   (nios_system_inst_sdram_wire_cas_n),                                      //                                   .cas_n
		.zs_cke_from_the_SDRAM                     (nios_system_inst_sdram_wire_cke),                                        //                                   .cke
		.zs_cs_n_from_the_SDRAM                    (nios_system_inst_sdram_wire_cs_n),                                       //                                   .cs_n
		.zs_dq_to_and_from_the_SDRAM               (nios_system_inst_sdram_wire_dq),                                         //                                   .dq
		.zs_dqm_from_the_SDRAM                     (nios_system_inst_sdram_wire_dqm),                                        //                                   .dqm
		.zs_ras_n_from_the_SDRAM                   (nios_system_inst_sdram_wire_ras_n),                                      //                                   .ras_n
		.zs_we_n_from_the_SDRAM                    (nios_system_inst_sdram_wire_we_n),                                       //                                   .we_n
		.GPIO_to_and_from_the_Expansion_JP5        (nios_system_inst_expansion_jp5_external_interface_export),               //   Expansion_JP5_external_interface.export
		.LEDG_from_the_Green_LEDs                  (nios_system_inst_green_leds_external_interface_export),                  //      Green_LEDs_external_interface.export
		.PS2_CLK_to_and_from_the_PS2_Port_Dual     (nios_system_inst_ps2_port_dual_external_interface_clk),                  //   PS2_Port_Dual_external_interface.CLK
		.PS2_DAT_to_and_from_the_PS2_Port_Dual     (nios_system_inst_ps2_port_dual_external_interface_dat),                  //                                   .DAT
		.Slider_Switches_external_interface_export (nios_system_inst_slider_switches_external_interface_bfm_conduit_export), // Slider_Switches_external_interface.export
		.I2C_SDAT_to_and_from_the_AV_Config        (nios_system_inst_av_config_external_interface_sdat),                     //       AV_Config_external_interface.SDAT
		.I2C_SCLK_from_the_AV_Config               (nios_system_inst_av_config_external_interface_sclk),                     //                                   .SCLK
		.PS2_CLK_to_and_from_the_PS2_Port          (nios_system_inst_ps2_port_external_interface_clk),                       //        PS2_Port_external_interface.CLK
		.PS2_DAT_to_and_from_the_PS2_Port          (nios_system_inst_ps2_port_external_interface_dat),                       //                                   .DAT
		.KEY_to_the_Pushbuttons                    (nios_system_inst_pushbuttons_external_interface_bfm_conduit_export),     //     Pushbuttons_external_interface.export
		.clk                                       (nios_system_inst_clk_clk_in_bfm_clk_clk),                                //                         clk_clk_in.clk
		.HEX0_from_the_HEX3_HEX0                   (nios_system_inst_hex3_hex0_external_interface_hex0),                     //       HEX3_HEX0_external_interface.HEX0
		.HEX1_from_the_HEX3_HEX0                   (nios_system_inst_hex3_hex0_external_interface_hex1),                     //                                   .HEX1
		.HEX2_from_the_HEX3_HEX0                   (nios_system_inst_hex3_hex0_external_interface_hex2),                     //                                   .HEX2
		.HEX3_from_the_HEX3_HEX0                   (nios_system_inst_hex3_hex0_external_interface_hex3),                     //                                   .HEX3
		.clk_27                                    (nios_system_inst_clk_27_clk_in_bfm_clk_clk),                             //                      clk_27_clk_in.clk
		.audio_clk                                 (),                                                                       //                              audio.clk
		.sdram_clk                                 (),                                                                       //                              sdram.clk
		.irda_TXD                                  (nios_system_inst_irda_txd),                                              //                               irda.TXD
		.irda_RXD                                  (nios_system_inst_irda_bfm_conduit_rxd),                                  //                                   .RXD
		.sdcard_b_SD_cmd                           (nios_system_inst_sdcard_b_sd_cmd),                                       //                             sdcard.b_SD_cmd
		.sdcard_b_SD_dat                           (nios_system_inst_sdcard_b_sd_dat),                                       //                                   .b_SD_dat
		.sdcard_b_SD_dat3                          (nios_system_inst_sdcard_b_sd_dat3),                                      //                                   .b_SD_dat3
		.sdcard_o_SD_clock                         (nios_system_inst_sdcard_o_sd_clock),                                     //                                   .o_SD_clock
		.flash_ADDR                                (nios_system_inst_flash_addr),                                            //                              flash.ADDR
		.flash_CE_N                                (nios_system_inst_flash_ce_n),                                            //                                   .CE_N
		.flash_OE_N                                (nios_system_inst_flash_oe_n),                                            //                                   .OE_N
		.flash_WE_N                                (nios_system_inst_flash_we_n),                                            //                                   .WE_N
		.flash_RST_N                               (nios_system_inst_flash_rst_n),                                           //                                   .RST_N
		.flash_DQ                                  (nios_system_inst_flash_dq),                                              //                                   .DQ
		.video_in_TD_CLK27                         (nios_system_inst_video_in_bfm_conduit_td_clk27),                         //                           video_in.TD_CLK27
		.video_in_TD_DATA                          (nios_system_inst_video_in_bfm_conduit_td_data),                          //                                   .TD_DATA
		.video_in_TD_HS                            (nios_system_inst_video_in_bfm_conduit_td_hs),                            //                                   .TD_HS
		.video_in_TD_VS                            (nios_system_inst_video_in_bfm_conduit_td_vs),                            //                                   .TD_VS
		.video_in_clk27_reset                      (nios_system_inst_video_in_bfm_conduit_clk27_reset),                      //                                   .clk27_reset
		.video_in_TD_RESET                         (nios_system_inst_video_in_td_reset),                                     //                                   .TD_RESET
		.video_in_overflow_flag                    (nios_system_inst_video_in_overflow_flag),                                //                                   .overflow_flag
		.camera_config_I2C_SDAT                    (nios_system_inst_camera_config_i2c_sdat),                                //                      camera_config.I2C_SDAT
		.camera_config_I2C_SCLK                    (nios_system_inst_camera_config_i2c_sclk),                                //                                   .I2C_SCLK
		.camera_config_exposure                    (nios_system_inst_camera_config_bfm_conduit_exposure),                    //                                   .exposure
		.camera_in_PIXEL_CLK                       (nios_system_inst_camera_in_bfm_conduit_pixel_clk),                       //                          camera_in.PIXEL_CLK
		.camera_in_LINE_VALID                      (nios_system_inst_camera_in_bfm_conduit_line_valid),                      //                                   .LINE_VALID
		.camera_in_FRAME_VALID                     (nios_system_inst_camera_in_bfm_conduit_frame_valid),                     //                                   .FRAME_VALID
		.camera_in_pixel_clk_reset                 (nios_system_inst_camera_in_bfm_conduit_pixel_clk_reset),                 //                                   .pixel_clk_reset
		.camera_in_PIXEL_DATA                      (nios_system_inst_camera_in_bfm_conduit_pixel_data),                      //                                   .PIXEL_DATA
		.lcd_controller_external_interface_CLK     (nios_system_inst_lcd_controller_external_interface_clk),                 //  lcd_controller_external_interface.CLK
		.lcd_controller_external_interface_HS      (nios_system_inst_lcd_controller_external_interface_hs),                  //                                   .HS
		.lcd_controller_external_interface_VS      (nios_system_inst_lcd_controller_external_interface_vs),                  //                                   .VS
		.lcd_controller_external_interface_DATA_EN (nios_system_inst_lcd_controller_external_interface_data_en),             //                                   .DATA_EN
		.lcd_controller_external_interface_R       (nios_system_inst_lcd_controller_external_interface_r),                   //                                   .R
		.lcd_controller_external_interface_G       (nios_system_inst_lcd_controller_external_interface_g),                   //                                   .G
		.lcd_controller_external_interface_B       (nios_system_inst_lcd_controller_external_interface_b),                   //                                   .B
		.vga_clk_out_clk_clk                       (),                                                                       //                    vga_clk_out_clk.clk
		.accelerometer_I2C_SDAT                    (nios_system_inst_accelerometer_i2c_sdat),                                //                      accelerometer.I2C_SDAT
		.accelerometer_I2C_SCLK                    (nios_system_inst_accelerometer_i2c_sclk),                                //                                   .I2C_SCLK
		.accelerometer_G_SENSOR_CS_N               (nios_system_inst_accelerometer_g_sensor_cs_n),                           //                                   .G_SENSOR_CS_N
		.accelerometer_G_SENSOR_INT                (nios_system_inst_accelerometer_bfm_conduit_g_sensor_int),                //                                   .G_SENSOR_INT
		.usb_INT1                                  (nios_system_inst_usb_bfm_conduit_int1),                                  //                                usb.INT1
		.usb_DATA                                  (nios_system_inst_usb_data),                                              //                                   .DATA
		.usb_RST_N                                 (nios_system_inst_usb_rst_n),                                             //                                   .RST_N
		.usb_ADDR                                  (nios_system_inst_usb_addr),                                              //                                   .ADDR
		.usb_CS_N                                  (nios_system_inst_usb_cs_n),                                              //                                   .CS_N
		.usb_RD_N                                  (nios_system_inst_usb_rd_n),                                              //                                   .RD_N
		.usb_WR_N                                  (nios_system_inst_usb_wr_n),                                              //                                   .WR_N
		.usb_INT0                                  (nios_system_inst_usb_bfm_conduit_int0),                                  //                                   .INT0
		.vga_controller_external_interface_CLK     (nios_system_inst_vga_controller_external_interface_clk),                 //  vga_controller_external_interface.CLK
		.vga_controller_external_interface_HS      (nios_system_inst_vga_controller_external_interface_hs),                  //                                   .HS
		.vga_controller_external_interface_VS      (nios_system_inst_vga_controller_external_interface_vs),                  //                                   .VS
		.vga_controller_external_interface_BLANK   (nios_system_inst_vga_controller_external_interface_blank),               //                                   .BLANK
		.vga_controller_external_interface_SYNC    (nios_system_inst_vga_controller_external_interface_sync),                //                                   .SYNC
		.vga_controller_external_interface_R       (nios_system_inst_vga_controller_external_interface_r),                   //                                   .R
		.vga_controller_external_interface_G       (nios_system_inst_vga_controller_external_interface_g),                   //                                   .G
		.vga_controller_external_interface_B       (nios_system_inst_vga_controller_external_interface_b),                   //                                   .B
		.enet_pcs_mac_tx_clk                       (nios_system_inst_enet_pcs_mac_tx_bfm_clk_clk),                           //                    enet_pcs_mac_tx.clk
		.enet_pcs_mac_rx_clk                       (nios_system_inst_enet_pcs_mac_rx_bfm_clk_clk),                           //                    enet_pcs_mac_rx.clk
		.enet_mac_status_set_10                    (nios_system_inst_enet_mac_status_bfm_conduit_set_10),                    //                    enet_mac_status.set_10
		.enet_mac_status_set_1000                  (nios_system_inst_enet_mac_status_bfm_conduit_set_1000),                  //                                   .set_1000
		.enet_mac_status_eth_mode                  (nios_system_inst_enet_mac_status_eth_mode),                              //                                   .eth_mode
		.enet_mac_status_ena_10                    (nios_system_inst_enet_mac_status_ena_10),                                //                                   .ena_10
		.enet_mac_rgmii_rgmii_in                   (nios_system_inst_enet_mac_rgmii_bfm_conduit_rgmii_in),                   //                     enet_mac_rgmii.rgmii_in
		.enet_mac_rgmii_rgmii_out                  (nios_system_inst_enet_mac_rgmii_rgmii_out),                              //                                   .rgmii_out
		.enet_mac_rgmii_rx_control                 (nios_system_inst_enet_mac_rgmii_bfm_conduit_rx_control),                 //                                   .rx_control
		.enet_mac_rgmii_tx_control                 (nios_system_inst_enet_mac_rgmii_tx_control),                             //                                   .tx_control
		.enet_mac_mdio_mdc                         (nios_system_inst_enet_mac_mdio_mdc),                                     //                      enet_mac_mdio.mdc
		.enet_mac_mdio_mdio_in                     (nios_system_inst_enet_mac_mdio_bfm_conduit_mdio_in),                     //                                   .mdio_in
		.enet_mac_mdio_mdio_out                    (nios_system_inst_enet_mac_mdio_mdio_out),                                //                                   .mdio_out
		.enet_mac_mdio_mdio_oen                    (nios_system_inst_enet_mac_mdio_mdio_oen),                                //                                   .mdio_oen
		.enet_mac_misc_xon_gen                     (nios_system_inst_enet_mac_misc_bfm_conduit_xon_gen),                     //                      enet_mac_misc.xon_gen
		.enet_mac_misc_xoff_gen                    (nios_system_inst_enet_mac_misc_bfm_conduit_xoff_gen),                    //                                   .xoff_gen
		.enet_mac_misc_magic_wakeup                (nios_system_inst_enet_mac_misc_magic_wakeup),                            //                                   .magic_wakeup
		.enet_mac_misc_magic_sleep_n               (nios_system_inst_enet_mac_misc_bfm_conduit_magic_sleep_n),               //                                   .magic_sleep_n
		.enet_mac_misc_ff_tx_crc_fwd               (nios_system_inst_enet_mac_misc_bfm_conduit_ff_tx_crc_fwd),               //                                   .ff_tx_crc_fwd
		.enet_mac_misc_ff_tx_septy                 (nios_system_inst_enet_mac_misc_ff_tx_septy),                             //                                   .ff_tx_septy
		.enet_mac_misc_tx_ff_uflow                 (nios_system_inst_enet_mac_misc_tx_ff_uflow),                             //                                   .tx_ff_uflow
		.enet_mac_misc_ff_tx_a_full                (nios_system_inst_enet_mac_misc_ff_tx_a_full),                            //                                   .ff_tx_a_full
		.enet_mac_misc_ff_tx_a_empty               (nios_system_inst_enet_mac_misc_ff_tx_a_empty),                           //                                   .ff_tx_a_empty
		.enet_mac_misc_rx_err_stat                 (nios_system_inst_enet_mac_misc_rx_err_stat),                             //                                   .rx_err_stat
		.enet_mac_misc_rx_frm_type                 (nios_system_inst_enet_mac_misc_rx_frm_type),                             //                                   .rx_frm_type
		.enet_mac_misc_ff_rx_dsav                  (nios_system_inst_enet_mac_misc_ff_rx_dsav),                              //                                   .ff_rx_dsav
		.enet_mac_misc_ff_rx_a_full                (nios_system_inst_enet_mac_misc_ff_rx_a_full),                            //                                   .ff_rx_a_full
		.enet_mac_misc_ff_rx_a_empty               (nios_system_inst_enet_mac_misc_ff_rx_a_empty)                            //                                   .ff_rx_a_empty
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_system_inst_clk_clk_in_bfm (
		.clk (nios_system_inst_clk_clk_in_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (27000000),
		.CLOCK_UNIT (1)
	) nios_system_inst_clk_27_clk_in_bfm (
		.clk (nios_system_inst_clk_27_clk_in_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_system_inst_enet_pcs_mac_tx_bfm (
		.clk (nios_system_inst_enet_pcs_mac_tx_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_system_inst_enet_pcs_mac_rx_bfm (
		.clk (nios_system_inst_enet_pcs_mac_rx_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) nios_system_inst_merged_resets_in_reset_bfm (
		.reset (nios_system_inst_merged_resets_in_reset_bfm_reset_reset), // reset.reset_n
		.clk   (nios_system_inst_clk_clk_in_bfm_clk_clk)                  //   clk.clk
	);

	altera_conduit_bfm nios_system_inst_hex7_hex4_external_interface_bfm (
		.sig_HEX4 (nios_system_inst_hex7_hex4_external_interface_hex4), // conduit.HEX4
		.sig_HEX5 (nios_system_inst_hex7_hex4_external_interface_hex5), //        .HEX5
		.sig_HEX6 (nios_system_inst_hex7_hex4_external_interface_hex6), //        .HEX6
		.sig_HEX7 (nios_system_inst_hex7_hex4_external_interface_hex7)  //        .HEX7
	);

	altera_conduit_bfm_0002 nios_system_inst_sram_external_interface_bfm (
		.sig_DQ   (nios_system_inst_sram_external_interface_dq),   // conduit.DQ
		.sig_ADDR (nios_system_inst_sram_external_interface_addr), //        .ADDR
		.sig_LB_N (nios_system_inst_sram_external_interface_lb_n), //        .LB_N
		.sig_UB_N (nios_system_inst_sram_external_interface_ub_n), //        .UB_N
		.sig_CE_N (nios_system_inst_sram_external_interface_ce_n), //        .CE_N
		.sig_OE_N (nios_system_inst_sram_external_interface_oe_n), //        .OE_N
		.sig_WE_N (nios_system_inst_sram_external_interface_we_n)  //        .WE_N
	);

	altera_conduit_bfm_0003 nios_system_inst_char_lcd_16x2_external_interface_bfm (
		.sig_DATA (nios_system_inst_char_lcd_16x2_external_interface_data), // conduit.DATA
		.sig_ON   (nios_system_inst_char_lcd_16x2_external_interface_on),   //        .ON
		.sig_BLON (nios_system_inst_char_lcd_16x2_external_interface_blon), //        .BLON
		.sig_EN   (nios_system_inst_char_lcd_16x2_external_interface_en),   //        .EN
		.sig_RS   (nios_system_inst_char_lcd_16x2_external_interface_rs),   //        .RS
		.sig_RW   (nios_system_inst_char_lcd_16x2_external_interface_rw)    //        .RW
	);

	altera_conduit_bfm_0004 nios_system_inst_serial_port_external_interface_bfm (
		.sig_RXD (nios_system_inst_serial_port_external_interface_bfm_conduit_rxd), // conduit.RXD
		.sig_TXD (nios_system_inst_serial_port_external_interface_txd)              //        .TXD
	);

	altera_conduit_bfm_0005 nios_system_inst_audio_external_interface_bfm (
		.sig_ADCDAT  (nios_system_inst_audio_external_interface_bfm_conduit_adcdat),  // conduit.ADCDAT
		.sig_ADCLRCK (nios_system_inst_audio_external_interface_bfm_conduit_adclrck), //        .ADCLRCK
		.sig_BCLK    (nios_system_inst_audio_external_interface_bfm_conduit_bclk),    //        .BCLK
		.sig_DACDAT  (nios_system_inst_audio_external_interface_dacdat),              //        .DACDAT
		.sig_DACLRCK (nios_system_inst_audio_external_interface_bfm_conduit_daclrck)  //        .DACLRCK
	);

	altera_conduit_bfm_0006 nios_system_inst_red_leds_external_interface_bfm (
		.sig_export (nios_system_inst_red_leds_external_interface_export)  // conduit.export
	);

	altera_conduit_bfm_0007 nios_system_inst_sdram_wire_bfm (
		.sig_addr  (nios_system_inst_sdram_wire_addr),  // conduit.addr
		.sig_ba    (nios_system_inst_sdram_wire_ba),    //        .ba
		.sig_cas_n (nios_system_inst_sdram_wire_cas_n), //        .cas_n
		.sig_cke   (nios_system_inst_sdram_wire_cke),   //        .cke
		.sig_cs_n  (nios_system_inst_sdram_wire_cs_n),  //        .cs_n
		.sig_dq    (nios_system_inst_sdram_wire_dq),    //        .dq
		.sig_dqm   (nios_system_inst_sdram_wire_dqm),   //        .dqm
		.sig_ras_n (nios_system_inst_sdram_wire_ras_n), //        .ras_n
		.sig_we_n  (nios_system_inst_sdram_wire_we_n)   //        .we_n
	);

	altera_conduit_bfm_0008 nios_system_inst_expansion_jp5_external_interface_bfm (
		.sig_export (nios_system_inst_expansion_jp5_external_interface_export)  // conduit.export
	);

	altera_conduit_bfm_0009 nios_system_inst_green_leds_external_interface_bfm (
		.sig_export (nios_system_inst_green_leds_external_interface_export)  // conduit.export
	);

	altera_conduit_bfm_0010 nios_system_inst_ps2_port_dual_external_interface_bfm (
		.sig_CLK (nios_system_inst_ps2_port_dual_external_interface_clk), // conduit.CLK
		.sig_DAT (nios_system_inst_ps2_port_dual_external_interface_dat)  //        .DAT
	);

	altera_conduit_bfm_0011 nios_system_inst_slider_switches_external_interface_bfm (
		.sig_export (nios_system_inst_slider_switches_external_interface_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0012 nios_system_inst_av_config_external_interface_bfm (
		.sig_SDAT (nios_system_inst_av_config_external_interface_sdat), // conduit.SDAT
		.sig_SCLK (nios_system_inst_av_config_external_interface_sclk)  //        .SCLK
	);

	altera_conduit_bfm_0010 nios_system_inst_ps2_port_external_interface_bfm (
		.sig_CLK (nios_system_inst_ps2_port_external_interface_clk), // conduit.CLK
		.sig_DAT (nios_system_inst_ps2_port_external_interface_dat)  //        .DAT
	);

	altera_conduit_bfm_0013 nios_system_inst_pushbuttons_external_interface_bfm (
		.sig_export (nios_system_inst_pushbuttons_external_interface_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0014 nios_system_inst_hex3_hex0_external_interface_bfm (
		.sig_HEX0 (nios_system_inst_hex3_hex0_external_interface_hex0), // conduit.HEX0
		.sig_HEX1 (nios_system_inst_hex3_hex0_external_interface_hex1), //        .HEX1
		.sig_HEX2 (nios_system_inst_hex3_hex0_external_interface_hex2), //        .HEX2
		.sig_HEX3 (nios_system_inst_hex3_hex0_external_interface_hex3)  //        .HEX3
	);

	altera_conduit_bfm_0015 nios_system_inst_irda_bfm (
		.sig_TXD (nios_system_inst_irda_txd),             // conduit.TXD
		.sig_RXD (nios_system_inst_irda_bfm_conduit_rxd)  //        .RXD
	);

	altera_conduit_bfm_0016 nios_system_inst_sdcard_bfm (
		.sig_b_SD_cmd   (nios_system_inst_sdcard_b_sd_cmd),   // conduit.b_SD_cmd
		.sig_b_SD_dat   (nios_system_inst_sdcard_b_sd_dat),   //        .b_SD_dat
		.sig_b_SD_dat3  (nios_system_inst_sdcard_b_sd_dat3),  //        .b_SD_dat3
		.sig_o_SD_clock (nios_system_inst_sdcard_o_sd_clock)  //        .o_SD_clock
	);

	altera_conduit_bfm_0017 nios_system_inst_flash_bfm (
		.sig_ADDR  (nios_system_inst_flash_addr),  // conduit.ADDR
		.sig_CE_N  (nios_system_inst_flash_ce_n),  //        .CE_N
		.sig_OE_N  (nios_system_inst_flash_oe_n),  //        .OE_N
		.sig_WE_N  (nios_system_inst_flash_we_n),  //        .WE_N
		.sig_RST_N (nios_system_inst_flash_rst_n), //        .RST_N
		.sig_DQ    (nios_system_inst_flash_dq)     //        .DQ
	);

	altera_conduit_bfm_0018 nios_system_inst_video_in_bfm (
		.sig_TD_CLK27      (nios_system_inst_video_in_bfm_conduit_td_clk27),    // conduit.TD_CLK27
		.sig_TD_DATA       (nios_system_inst_video_in_bfm_conduit_td_data),     //        .TD_DATA
		.sig_TD_HS         (nios_system_inst_video_in_bfm_conduit_td_hs),       //        .TD_HS
		.sig_TD_VS         (nios_system_inst_video_in_bfm_conduit_td_vs),       //        .TD_VS
		.sig_clk27_reset   (nios_system_inst_video_in_bfm_conduit_clk27_reset), //        .clk27_reset
		.sig_TD_RESET      (nios_system_inst_video_in_td_reset),                //        .TD_RESET
		.sig_overflow_flag (nios_system_inst_video_in_overflow_flag)            //        .overflow_flag
	);

	altera_conduit_bfm_0019 nios_system_inst_camera_config_bfm (
		.sig_I2C_SDAT (nios_system_inst_camera_config_i2c_sdat),             // conduit.I2C_SDAT
		.sig_I2C_SCLK (nios_system_inst_camera_config_i2c_sclk),             //        .I2C_SCLK
		.sig_exposure (nios_system_inst_camera_config_bfm_conduit_exposure)  //        .exposure
	);

	altera_conduit_bfm_0020 nios_system_inst_camera_in_bfm (
		.sig_PIXEL_CLK       (nios_system_inst_camera_in_bfm_conduit_pixel_clk),       // conduit.PIXEL_CLK
		.sig_LINE_VALID      (nios_system_inst_camera_in_bfm_conduit_line_valid),      //        .LINE_VALID
		.sig_FRAME_VALID     (nios_system_inst_camera_in_bfm_conduit_frame_valid),     //        .FRAME_VALID
		.sig_pixel_clk_reset (nios_system_inst_camera_in_bfm_conduit_pixel_clk_reset), //        .pixel_clk_reset
		.sig_PIXEL_DATA      (nios_system_inst_camera_in_bfm_conduit_pixel_data)       //        .PIXEL_DATA
	);

	altera_conduit_bfm_0021 nios_system_inst_lcd_controller_external_interface_bfm (
		.sig_CLK     (nios_system_inst_lcd_controller_external_interface_clk),     // conduit.CLK
		.sig_HS      (nios_system_inst_lcd_controller_external_interface_hs),      //        .HS
		.sig_VS      (nios_system_inst_lcd_controller_external_interface_vs),      //        .VS
		.sig_DATA_EN (nios_system_inst_lcd_controller_external_interface_data_en), //        .DATA_EN
		.sig_R       (nios_system_inst_lcd_controller_external_interface_r),       //        .R
		.sig_G       (nios_system_inst_lcd_controller_external_interface_g),       //        .G
		.sig_B       (nios_system_inst_lcd_controller_external_interface_b)        //        .B
	);

	altera_conduit_bfm_0022 nios_system_inst_accelerometer_bfm (
		.sig_I2C_SDAT      (nios_system_inst_accelerometer_i2c_sdat),                 // conduit.I2C_SDAT
		.sig_I2C_SCLK      (nios_system_inst_accelerometer_i2c_sclk),                 //        .I2C_SCLK
		.sig_G_SENSOR_CS_N (nios_system_inst_accelerometer_g_sensor_cs_n),            //        .G_SENSOR_CS_N
		.sig_G_SENSOR_INT  (nios_system_inst_accelerometer_bfm_conduit_g_sensor_int)  //        .G_SENSOR_INT
	);

	altera_conduit_bfm_0023 nios_system_inst_usb_bfm (
		.sig_INT1  (nios_system_inst_usb_bfm_conduit_int1), // conduit.INT1
		.sig_DATA  (nios_system_inst_usb_data),             //        .DATA
		.sig_RST_N (nios_system_inst_usb_rst_n),            //        .RST_N
		.sig_ADDR  (nios_system_inst_usb_addr),             //        .ADDR
		.sig_CS_N  (nios_system_inst_usb_cs_n),             //        .CS_N
		.sig_RD_N  (nios_system_inst_usb_rd_n),             //        .RD_N
		.sig_WR_N  (nios_system_inst_usb_wr_n),             //        .WR_N
		.sig_INT0  (nios_system_inst_usb_bfm_conduit_int0)  //        .INT0
	);

	altera_conduit_bfm_0024 nios_system_inst_vga_controller_external_interface_bfm (
		.sig_CLK   (nios_system_inst_vga_controller_external_interface_clk),   // conduit.CLK
		.sig_HS    (nios_system_inst_vga_controller_external_interface_hs),    //        .HS
		.sig_VS    (nios_system_inst_vga_controller_external_interface_vs),    //        .VS
		.sig_BLANK (nios_system_inst_vga_controller_external_interface_blank), //        .BLANK
		.sig_SYNC  (nios_system_inst_vga_controller_external_interface_sync),  //        .SYNC
		.sig_R     (nios_system_inst_vga_controller_external_interface_r),     //        .R
		.sig_G     (nios_system_inst_vga_controller_external_interface_g),     //        .G
		.sig_B     (nios_system_inst_vga_controller_external_interface_b)      //        .B
	);

	altera_conduit_bfm_0025 nios_system_inst_enet_mac_status_bfm (
		.sig_set_10   (nios_system_inst_enet_mac_status_bfm_conduit_set_10),   // conduit.set_10
		.sig_set_1000 (nios_system_inst_enet_mac_status_bfm_conduit_set_1000), //        .set_1000
		.sig_eth_mode (nios_system_inst_enet_mac_status_eth_mode),             //        .eth_mode
		.sig_ena_10   (nios_system_inst_enet_mac_status_ena_10)                //        .ena_10
	);

	altera_conduit_bfm_0026 nios_system_inst_enet_mac_rgmii_bfm (
		.sig_rgmii_in   (nios_system_inst_enet_mac_rgmii_bfm_conduit_rgmii_in),   // conduit.rgmii_in
		.sig_rgmii_out  (nios_system_inst_enet_mac_rgmii_rgmii_out),              //        .rgmii_out
		.sig_rx_control (nios_system_inst_enet_mac_rgmii_bfm_conduit_rx_control), //        .rx_control
		.sig_tx_control (nios_system_inst_enet_mac_rgmii_tx_control)              //        .tx_control
	);

	altera_conduit_bfm_0027 nios_system_inst_enet_mac_mdio_bfm (
		.sig_mdc      (nios_system_inst_enet_mac_mdio_mdc),                 // conduit.mdc
		.sig_mdio_in  (nios_system_inst_enet_mac_mdio_bfm_conduit_mdio_in), //        .mdio_in
		.sig_mdio_out (nios_system_inst_enet_mac_mdio_mdio_out),            //        .mdio_out
		.sig_mdio_oen (nios_system_inst_enet_mac_mdio_mdio_oen)             //        .mdio_oen
	);

	altera_conduit_bfm_0028 nios_system_inst_enet_mac_misc_bfm (
		.sig_xon_gen       (nios_system_inst_enet_mac_misc_bfm_conduit_xon_gen),       // conduit.xon_gen
		.sig_xoff_gen      (nios_system_inst_enet_mac_misc_bfm_conduit_xoff_gen),      //        .xoff_gen
		.sig_magic_wakeup  (nios_system_inst_enet_mac_misc_magic_wakeup),              //        .magic_wakeup
		.sig_magic_sleep_n (nios_system_inst_enet_mac_misc_bfm_conduit_magic_sleep_n), //        .magic_sleep_n
		.sig_ff_tx_crc_fwd (nios_system_inst_enet_mac_misc_bfm_conduit_ff_tx_crc_fwd), //        .ff_tx_crc_fwd
		.sig_ff_tx_septy   (nios_system_inst_enet_mac_misc_ff_tx_septy),               //        .ff_tx_septy
		.sig_tx_ff_uflow   (nios_system_inst_enet_mac_misc_tx_ff_uflow),               //        .tx_ff_uflow
		.sig_ff_tx_a_full  (nios_system_inst_enet_mac_misc_ff_tx_a_full),              //        .ff_tx_a_full
		.sig_ff_tx_a_empty (nios_system_inst_enet_mac_misc_ff_tx_a_empty),             //        .ff_tx_a_empty
		.sig_rx_err_stat   (nios_system_inst_enet_mac_misc_rx_err_stat),               //        .rx_err_stat
		.sig_rx_frm_type   (nios_system_inst_enet_mac_misc_rx_frm_type),               //        .rx_frm_type
		.sig_ff_rx_dsav    (nios_system_inst_enet_mac_misc_ff_rx_dsav),                //        .ff_rx_dsav
		.sig_ff_rx_a_full  (nios_system_inst_enet_mac_misc_ff_rx_a_full),              //        .ff_rx_a_full
		.sig_ff_rx_a_empty (nios_system_inst_enet_mac_misc_ff_rx_a_empty)              //        .ff_rx_a_empty
	);

endmodule
