// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
mH8NaBrdgAQDwF8FemNWZS424pk/zGPmBIi9YVjQvAHb+uPTKEaJNHjRlI5c/piphckTqvHo2MNM
yAkpuCKBgQ+sYjNLAtMFwt+8gfgewQngVUeDAOBpsDQkoz1G2bIzjg4C+RWkwswXKmRs2/sL9exl
+T/JJ27Zzwyu5eH4OnI7tXqWbPHW0VAkXj1nn0DRIDCBuW2IcO1cwf9ObtDV36LMVyrQXJfIGmKx
QawGa/5D2L1KHsOEAcIQ2xJtBBeAIhuycgSLG+MVs/WxzFgEPGnhtamM0ySKrbhdjy73aW9yn2eS
n/9tMomfCnHhkfFgyCOrjKJSnNGoHRGwJTjzGA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
rrKfBz2jrMr2lRIaavgfcd38ZMPIa6vzOVS5hd0uXFx7CnAZ+czFBQ+HoFDeU0qOqKSfGFVyhVDq
T77qFfKPMKqnUNVyJ1Ucb9UZgUdeaGquErEXV8G5VzkxghLNOQJ2A8Axe2EqeCm0pSX9CKnnALko
mzjidIBhMRrd0rx1Sqhfn6IZq7lrp9YSjJ4S7UFaLdxD/kJtAtN71RreHFs4UeUQFoRhaXTyRpdc
N6MBESbMqvlVy1Qzt4ETzf90//OmKueQktk1r1ZY8lS/AIDHRrWzJFjRgsuOfrU8jrWJGWJTYz6P
mhOeHSztxT2e0ayaJtmoRnGa+vaXcgcg5zhgI/Qc67Tdy3KDo8XWWh2EGAIq3fafMnbtcq5Pk4PF
nCJTpmgKAGUEnEddaX+fpvaW1rvOmrtr2uFVL7+vRl7D42xbilYUH+nu8Qu4iNVzekPR3yWZw38E
htjnzRtQh1kH0QkHhC1bSB3pt3y2l4FjTj5Ut1yt5q7mRC1hN6HJhrW+rMG2njBZHrfSsuF7JQH1
UZoeYT+GVSVAFHuEsvZK0DAn24o2nQq0VHol844Kc+BarVRh6a/UU46Eb4yXSr3C+OWRwJTiBsl+
AO+slFAZjmq1objAgSdaODH39NRtPUkfK92u/t93MqcRpaIzrCVoVgWls2wAiWaWPUclukcHH/GW
uQNoqu1bIT++jrrl0CFpycX1IxuZjmVTtxxtB0m/OTLSZcVogro/lIACvW21pL5YQnZCl/kY0KK0
UdmSNRbd7HHCF5yboUGjba1mzlCztZ1C2+iLqd9fxybEQwcIH+LQ/c3qdwEeMD9oFVW/1UAv1L1U
W+uqUlEr7swDDEAz/HRJQTve8t5moB0UQttbvx1xhCJAOc36q3EZwJor0EIjHSRX51WNN0Y4eQbj
ZcLYPvNt0vkLFJmMBQB9GROvqyaY2pnhWzWShmo9p/b8TsMcebdE9ji/PgyFZFWuUKHBstHgHil7
W+zmDbCmt3+RSlJuIAzCFb4TlBLBRq3d2r0M2t+tbnYEcGEcAU++9L1gy0jLChJ805St5j7EQLwg
tG8zwuRrDc5768l63Bz7UbkiWN4gJrD3z7QIE8stAE5/W1ib7c2fH5BSILDYv/0Hdq0LmDYaQXZG
qbM8/vUklwMztpKNAb1xsglZoOsQHiL1sCxKpkFs3e7pGsnWDhb6joLgDE8GznGBzzlckMelbaLw
4GhkPSlnVhv3bJGKai04lxUNHAz/krBi181YEV/hMn7wKpa60CluIb2+WTfJSTungyaLHsr6Pd4w
7MWFZLlKu/kdD1SBWf+22wkcek1L0eSc1GMAB/XhUGIbHtsdAcm30NcidyP/t4eIvQE3g6EdUIC6
hV7N8yVYbPOopxaLt7jDnHCUIRs5nv/ttON7Feo4OM7+vsOlHlSWHgOmwoTplxL7tofSUQ/CUtUe
fsfcZrYg+x/PPZc9sdnicf0iiieVzJhfzOMQifLWu29bdbJZjeHhYoRojM59tXmSNsGuOCi8kcYi
6cm/CV78iiAW3qqEMJK4b9gvLKwC5+SLsg02JwNdttyBkK8cEjTMr1+Q4qiE297NqtKQ8QPZ7Vxt
xVznacx3Txpe79uRf6EoSAideQ6mBkQFBQx2XtWTRv4GZxEAiiHMlbchYfgJdpbDdLLxtl257fbW
UyA8QyRMIS0dX6nzSXEoPG7UPnkBD0hMMGB3IeSLxUZdc+dqDCHApi8/cNoHyC4dZXXf9pvjL6G9
3JrrgmKNBkAJGUNqfe+0Q3eUvaMcG5oY7nuMHwyWAlU75MNactU1Va8WOBIK5Iu5sEm0/vX0OUWv
fW2IC0+UnaofrSobAgHzHyKdsbqeyct7P/4P7BY8B1BlE/Urm4rm4djdmrYUEOjx1bsXENdevevP
e/e+ciN6Xcb1M2eu9OTXwAedqwSQWOzl2fHP0iyCXe2dMryMu+NlwOCp2I29klNL49R3x42bl9pv
ZWDMgCl/ntZIF6MoGL+RmJwQtaLjDRJtEhJA6RxzhutrLwRRbMR5h9uXHWmFiMG9LZMEebsoS5VD
pM3iZy5Sp6h04ZOIenO823NZoMbDZs4HRXFsfns4+Jgd/oOy3S9WWYPyXzfNGF8IHGdyDWIW/cCE
VQt8yDrCk9sclOrblWiJ5HBq0hHPnDSu25vUF22QWAeHR/NZgafrs/tBpPYXahTIlMI8fw5LGQXO
Vnc/tgajQyL96uYiii7lBJqIf4UwAavKpYKZeLbYIaeB8o6vLzhk1A93syOkNR4jnjj+0KnTE7pp
R/ceIkVu+Z8ALoNubF746fwYKhuYekJQHiwFSP+ARdYq/VDt2irkwThE5qwMhVqp070NMzc5/XM3
W25p4vx1hIDALAiMqAx3ZFaCme58jL/NlHAGooPno2Pqb5YQ8G8IsWLjI0SdUJdhtvrQMSRxF3Yr
f2rBRaddlbTuc1EfV51Tl6kAc/hAYNbrePUs03vUkaErT3oXqHcSCRM7nCizHXOxREq5RnAan1sI
wTyXvTY4iJNtLQ0G2KJn75g6oYcXbTCycsoWrjPmtWt6IVvOtOl09GTWC7htITBTFQKLbiC0waf6
TreRRQ7X7hU6yoWrAHqK1rU58UDW+Z6Imq8J517rpYEYsdmH7XduNNAWKamVZUKoL1SNu1+6Zifd
xZuczT0F5OhY3ibNiNs82EQwicUU8v8TL4IVRIEW6F8Unp69yv7hnrAv3GSjWPDY217mcad3nhd7
+H4SRsCkkT3X3RZ/XRwaWjWbQe4G8LTo32OtgSzBAsdQ9mfIGaEImB+T2WdqKjxyJNEjg1dN0GjF
CnV9cduCcjey34svyOoKcskz4pFiqY/XLnVyZn9xYj7kr9H1YPnFQmEcF6tGFhmWsr6kVDcQ/m8G
e2PsgmOHDf0b30GC+CAVYRDGd/7bsPjI4oxNPTEqW/jU+4jHP4cL1grMKhQGpAKxhApkAQlJWD97
IYublKKppY+d5b5ZY2Xa4t1C/YDz2/hSL4TTI6zAg70uUc3K5Wvn0vvSDJ46+CPuPuf9zAEN34AX
ME4ISoqGkkyW9wRXWGdUlNg+C/LXuNnwS0d7v4AA4wsX6oIxUg7vmFlobrTSBoHhXP7wWyPmYs8l
6UOZcRu6yq5iyEnhI6z9sfsBYLSVcnf+F84qWVOVsmKWFwuj2MgfKVHxgZ9aVJ4+QYQ2i2rt3Y/r
TyKftQQw9UQWSXNtCUweJaSM5g8Gd7+MPTY8cF1uwVcgVWaGRQFLC9wPx1WlpObHmnZFf9Tg509f
OIm+I2FHFo61oWWDAqkRZDPSoMpfDsTMqdEQLu9Lo3wBQQi36kJ+adwYJ7bQka3Zn4uYf5Ds9kce
2csf/Bs6aao85s+oxrsH30FyRqL1pahrx/eEfZ5mkZ5SvkrFetVb6var3FB0Uvk6GVYFxGu83287
PkklH/B9TKRb9coSI/ec/gtyafyqDu/v0j24qVSB7BG4BtWexz4ywPP8WERmcfTr7q/l+eyrZz9Z
W1qf4JeMESDh4OF/InFeki8PY7EUQNEU7gsfhokH0IJSTifM8IdTFuoAEUy5H90XDcL25doIXN+S
BF5GfgWXdFYE89WzGpmg0oIXD5tg0Wj/KRX67LB45ZlnlfsQ8NfY3jbpuvE+AEcZpJYuDe6rWHRa
do6qHuaw9wmfTdHv5OatZ9qfPOpfJpPKkM7jXg0LzfIkplI1rFj/Q/DhHWx2bxwWOC6LculWII9v
irhAc6ZrDREWvfam2lHvMHgJKQ5XgGczlRenMmcmNp0eGuItvvWXvdZ11decXxFXRCN3AwEh9Vba
PIEExh1mlrlE8Wyc7b9tqq46jnRBX6Ttc5+OnKCLvPtDK9wlPBt+R3WzDkjYWtqdyS7HATEJZYY0
o8r7I0zRf/MVINF9CFUEyEZUTeJe8x7gAHTfUXexqdB74OyX7A4HighmSr53Msr+8HVqbB5QwbS7
gc5dGvEE/ewqTTa0EOhbLK0dW2qpB6/vJsyrFN6AIpwkvYJWU6bV92rwpJo4p7qPJJ2LcdTZ2DdI
F+c2CYP9wm7z26lotr0yy0f5CEqggrJiMvHpbSGBDWMgzuKTUTW3gxBD1/ZU4TN1n6cvWAnU0+5/
N15XOKSH8bPGs5HUk31XVk7nxSbmveH5xiyaomEn7K6sJjsTGrzkZFiWWeq/MByTQuFJfpFAd5Ua
i8Gwixx+liZEDm7B4jZzUYCLdbLlsQ48t4FtGevGbvhr4rFpaMaiM+nB7E14z95HNkqfFsIqE7QK
PusUJiSeqNR9B3ieYk6TWYLUcZPIkxEHc5JKrxikWLo/+RADkNkQAPnZd/zthhwbYJa/lbOSeLPu
1qIzRt/CDFGnMWX+HWLlmruxOWxo7Ie3hOc5mOFPuIS3uYKx1WrOHLiXoebxEZtRrBG2h9jOmLwU
6X7aQcJC/oUYZBakpn5Q1tTqY3OInRwGlbT9We4ORBNa744t9sm8NPTaD9uyQb3QrjNJ0mrUo/Gz
q1o0izzOWtA8POQhP/+eToPNCBkuMHWqStOEYcyYYJcf0qQwUxJl2RK+KCAMvo4hjPIDrRe/yB7Q
haXk38GqzM7XIvtJk50MVde5RH+fuBNFGr4d8/UbASSfPJlqpLXk/ZqmqtOCsWgptjncU5dw3M2M
T5hKTYwmKN6LsyR0c31VO98VkTxgi93mW3ygohlRrdGbyLTkC47OsjweJWkHEErW6AvRLIByFniu
1HdgULJUnYCbswkkPjErMjrUXIqcqtHI6SPDorOTAuUDf0iZitqYc52FKP4qGXJR57mPoGuxxxqF
Wi3uBu6zzC4lqIzNZ02vwZkjH1mOzEErG+9qvtP7EWGEP+aj6TQLKC+cPiILMjsqmG36A4yzIDE6
/iJyQfeDJ2YvlFM8GhEZSaSZMF7wXrokx+ja09MIkRLyVTya1KBPyCHIEktqvIVhiMi2iFn1mXZV
f925Mr58JFRcEXqZrl6AV9y6Kt/We0SrfxiFcaPS1uy1OBEREC5mxCGZeItTT/qI0YpsIEDw+fhu
M4qkxsciqzDYdoQJi4RA/1NUqu8BZEQjDOgcTDNw+VWREO3Dd8HcsGuZj4/bgL9UgM3rKGyE5l9n
ISKo8IIlINe3db3ITDs1wIKmh3s1kGCSaxG6hoWT4o5HtdBHxsFc1tajCKXCbL3j5WNP5JYcQ5On
J2Q1/DrVXTOtLsPWLsrLcse5Jo/KmTh6BBsjNp1+KH57/TQmiPHG3P+y6+mi3Z+bDubclZ0c9kTI
FRRAuKUQk3mDCf2Qsx6i2YywIU+syip/ZgsCDS/VWSEmVif8BsI7NwFVcScfk95ccEYqziIhjBa0
qJpm0l1GKX7QedLbUpL/Qd8HTwbg95AMPz1MFUvzD46rB4W7eaOma3AH9cR4rELVk5ty/6S5e++W
T/Ai2ganh03PWGNIgnVPaSSyVx6osb8izL2Bsfz9DSWLHmee+GvyNQR3u+EMOS3WFoCnvfY3DWot
odoaiNRUun3a4Tr7A69q2Twk6js09X/wqc7iJTNPsPFAvuh1FbAw5YiKu/cquQk/rewXqV8Kf8VD
lKmbpND+l5SGPJkkJkwskVDlEo9V/kFw0HsJeq5d/NhoeCqUTtiTK0KMHsEQ4/+oEsWsETTsJ97F
/LdZXRDnp3f0rAoyvDPJXdUj/SjCAAKONvKlJX4SVgiVUcsggeqF/TeI/D7FiF1dVDFBpfNCmmXL
gYxzAcBE3fhGCVWIqjT7ygpLGzzU7XxyZX1sKu2X8kjPFIvn8l/bEhatPciLXVvRuGAxaxL1YMdW
0Rkm7FkY50Ov5PkduoHCbKc0jMJycsveiB612jMxj2HWCgRM1AvYYsh3R5h2ojMdDluHoqcE+UOp
ycJ+gYdlemeKR+jKfraFW5fX+qGySxxa5aQIgYTweGDOeJF6l7pRpnQP94eR1YjHtCS9Wk14OUsx
7Bnr5Bxa5/epQI4gXr0UttFRLoSrfkWz2lZSSSJSNV43bqB9LI9fRXAy4MC/NBja2ST5taJ5DgN6
29F1ffoyFE3n9z6sdezE6z9NFnLtuIMsjSIXfQlnFp9+IvcWzFKjtBU/TcgEp8KSm6KZ/mNrJ8FD
0PaNCPeO8seId5ami78Ofmxy1O1i+6f3A3cFbcdRi5NjK0+K2qInOGDpJS2aA4ZTuyNt2w7lK5kT
gynnk9x3iSsS/UDLpnSgrvBj5l+2NYEJBWzeCVoMvzEOticV/76kQUeSxEYW1QsbxCXMnazVcwwN
fnij5bq/f2RHiGg5nLoyxXiHMrllqq4zoKrQd0txKv6FZgQGH3zfNYSLRrU/9zbEAi74DcOQa74H
Z/75knpIur9z1EOZGsCgjyfSDCyaX3/G+l8+NLtueNDKxfoRRskpPPYrwc3rF2kaTNE9K57yk2Tz
4RV5sy2rAHmVaLDkFiVfgbrclOcwlSNSPY1/cgvB40rVAdx+QsCb+7sa+vUgoKZuX9od+2w9PuvK
v59jSn66aTbWVLY3wH35KrXnc8BN5MNSoxEe8Z4xW0jIkAV6BSsvSDNrO9lJ/a5IPXydIyCIAHg6
1BEFYk9r46CtuawewTcp8XJPWbfIQ5byC4FHrJVBGbGIkRhzd3/FBcQfsn6eUqVcbNaT55h+y8RU
mJQpxEIQod8BdMpORac5KPKTGK28q4viGzEdcHin25JidDUc7vq2AyUyxkEtpNEwSyWWyBeixHDq
eviJ5fuxjjiXiko/RegLsv+AEhAIisBNSPB5ty36uCKhH3XGOgi2p61rD9FHbgFxDoC15hVOOuKx
DXak8w8u9FoEwPJ9XZW+aYvCWLtD6P43JG7UVHNsOawRrkL7kvM2TXRA7P5rabWb5J2QaAeWEGLe
QHvlIb8XWzYN1MbGCTTou4fEZFPmKZcRfoKJy/oZYCwsGQjiYBh7SOpBSx5SZzOP5CRPsS6dp5m3
DL8g7E0OS8mWaylAO5rsrnrSmFUiiLPe71DnY5uwr9N5p9ca4h8k6H+0T6iCrwvK5W4n+OA5R5Ok
w801egnTvCkmchdyPByGHppbIqTZdvJazPNSTodNZ+0P1cqejxoKlSTFxDXblhDZVgFs6ASexfbp
e7KEz0ipLrboIZrl+55FBPXBRU24mVSvjX2l4hM/25mjTVctik4jtrVi3YPpiVkuTV4um/rVnG74
1EY7Xh5UJMW2syd47YvsBQbiIylKBJhK7uBma/AhD2IukB8xacSwFkPt3HWY4z1zexhw1NCve+Or
DDQrd6jYgpaNXgcJ0gTIni7BxytJwbEdw2q1SdJfmi8Ap1bzpEzCF6DBnQnPr5ybDq2vPSyHU8g4
clc06nPeY4IwsP563sVibaIL0A112YbnHiBAZkvcqkam/c29hDxT/x5GKFCqSfTSD9Odcoemk/Ei
PAACyaA5BQKeo3/Qf/zrHW/ngL2rgdVHkS04Tl5a0HnkQy60i//N7urpoEo5357v13gTd6gFT7Oe
Uprx1/1u3IU2UqPDpfhirgpe1sSkAjZnUEpuoevaFM6LKcqVRn1HbcssFal0+2FSLdZvF/NDlKGD
nZRohVo2rWrDupnrCeI9+JTQHmzUjU4UUvXfkWx5SmmDWjD4V2w4x5Jo+IXBPvqCqi5Dru7ZqTuI
Xl6HvgDMW7plakZa8hbhgiU2HMDyiwR5kHFT2DklkAcr0gJZn1ZTeNO9V6xXNq45WYsbfXdVMfzt
yxdcrSdUV3xvNsDk1KLI/Uu+J5RXbWgkbwXMzsnt3Mi2O7zQQ5DSrNOH61nET0QS9XKdTAdiVssV
MU5iHCjVamWqUtJBDC6UIO0f624IKpGoUoe0Lwy9cWebAfb3Vq1j7M3iZvwAnYJATCre8O1WY1N0
QTQCSm9YIylDkDSM9StIIfRi15MucLNfNe4bctB9OBqGtq2h3k+Wvcf8aruT2PfLjtq8TS4kXvw0
MN7Ng+P0g6xY2ck8X5b95U5flHoLUkPm3k3XLYtGDn6ejrfc2FJs7htddd1jBQYKEODzgF2Lsrys
6Tz3FCGwANbVFx50we+ol9OUxZXwqLiwD+/GG1Xh7oOioMIiuSOSFmicOxXL72rF+VblHL2tKhIl
RNdNUS3c3N1M9L/pU3HLr6aK8N9LeClbChksOclUQfM8D1PzytL3mQFywURUulAddIOnfzGsjugr
mPhi4S4iq14CAS6nywrXb7jEESgylprHPtD0Wepvr6EQ5C9s2UCBCLCGLnNakztbgPuiSy/9Bced
KW8k/v8l0JcmRwiiB44H7Bme7wAaakVmC/zxUcHlmOXMbuvZRKlYqJyzpsQ/46euFVhhwlbtnRm0
AsGulXrz/9hqkYx+PXczj7VtouQrCM9CYkQy/yLoPpCs2NfxHMEbToQ46QUUQXIx7NTKqO8gbCL4
HoZw2Obkg/kIQLffZ7xugMVB0NSJF2of9cDpfE9RrRrOVlciYOPk8N2GMdogAcGoiwRmW8AjLdaX
aVisbinz5Vkd
`pragma protect end_protected
